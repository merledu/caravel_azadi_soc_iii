##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Tue Mar 22 08:11:57 2022
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2299.540000 BY 2118.880000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 345.514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1843.68 LAYER met3  ;
    ANTENNAGATEAREA 0.852 LAYER met3  ;
    ANTENNAMAXAREACAR 406.125 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2165.77 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 6.380000 0.000000 6.520000 0.485000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.771 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 151.239 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 755.223 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 4.090000 0.000000 4.230000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.050000 0.000000 471.190000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.320000 0.000000 158.460000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.625000 0.000000 475.765000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.475000 0.000000 466.615000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.795000 0.000000 461.935000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.220000 0.000000 457.360000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.160000 0.000000 453.300000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.505000 0.000000 303.645000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.825000 0.000000 298.965000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.250000 0.000000 294.390000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.675000 0.000000 289.815000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.100000 0.000000 285.240000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.420000 0.000000 280.560000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.840000 0.000000 275.980000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.785000 0.000000 271.925000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.105000 0.000000 267.245000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.530000 0.000000 262.670000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.955000 0.000000 258.095000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.480000 0.000000 253.620000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.905000 0.000000 249.045000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.225000 0.000000 244.365000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.650000 0.000000 239.790000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.595000 0.000000 235.735000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.020000 0.000000 231.160000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.340000 0.000000 226.480000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.760000 0.000000 221.900000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.185000 0.000000 217.325000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.505000 0.000000 212.645000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.930000 0.000000 208.070000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.355000 0.000000 203.495000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.195000 0.000000 199.335000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.720000 0.000000 194.860000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.940000 0.000000 190.080000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.465000 0.000000 185.605000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.890000 0.000000 181.030000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.315000 0.000000 176.455000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.635000 0.000000 171.775000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.060000 0.000000 167.200000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.000000 0.000000 163.140000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.745000 0.000000 153.885000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.170000 0.000000 149.310000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.595000 0.000000 144.735000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.120000 0.000000 140.260000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.340000 0.000000 135.480000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.865000 0.000000 131.005000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.705000 0.000000 126.845000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.130000 0.000000 122.270000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.450000 0.000000 117.590000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.875000 0.000000 113.015000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.300000 0.000000 108.440000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.720000 0.000000 103.860000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.145000 0.000000 99.285000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.465000 0.000000 94.605000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.410000 0.000000 90.550000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.835000 0.000000 85.975000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.360000 0.000000 81.500000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.580000 0.000000 76.720000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.105000 0.000000 72.245000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.530000 0.000000 67.670000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.850000 0.000000 62.990000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.275000 0.000000 58.415000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.220000 0.000000 54.360000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.540000 0.000000 49.680000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.960000 0.000000 45.100000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.385000 0.000000 40.525000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.810000 0.000000 35.950000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.235000 0.000000 31.375000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.555000 0.000000 26.695000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.980000 0.000000 22.120000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.820000 0.000000 17.960000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.345000 0.000000 13.485000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 8.560000 0.000000 8.700000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 448.480000 0.000000 448.620000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.973 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 443.905000 0.000000 444.045000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 439.435000 0.000000 439.575000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 434.860000 0.000000 435.000000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.721 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 430.180000 0.000000 430.320000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1792 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 425.600000 0.000000 425.740000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 421.025000 0.000000 421.165000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 416.865000 0.000000 417.005000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 412.290000 0.000000 412.430000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 407.715000 0.000000 407.855000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 403.140000 0.000000 403.280000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 398.560000 0.000000 398.700000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.749 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 393.880000 0.000000 394.020000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 389.305000 0.000000 389.445000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 384.835000 0.000000 384.975000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 380.675000 0.000000 380.815000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.84 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 375.890000 0.000000 376.030000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 371.420000 0.000000 371.560000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 366.840000 0.000000 366.980000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 362.265000 0.000000 362.405000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.854 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 357.690000 0.000000 357.830000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.798 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 353.010000 0.000000 353.150000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 348.435000 0.000000 348.575000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 344.380000 0.000000 344.520000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 339.700000 0.000000 339.840000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.833 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 335.120000 0.000000 335.260000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 330.545000 0.000000 330.685000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 326.075000 0.000000 326.215000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.214 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 321.290000 0.000000 321.430000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.214 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 316.820000 0.000000 316.960000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 312.240000 0.000000 312.380000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 308.080000 0.000000 308.220000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.945000 0.000000 1056.085000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.475000 0.000000 1051.615000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.900000 0.000000 1047.040000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.530000 0.000000 1042.670000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.060000 0.000000 1038.200000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.480000 0.000000 1033.620000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.905000 0.000000 1029.045000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.225000 0.000000 1024.365000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.650000 0.000000 1019.790000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.075000 0.000000 1015.215000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.500000 0.000000 1010.640000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.920000 0.000000 1006.060000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.760000 0.000000 1001.900000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.185000 0.000000 997.325000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.715000 0.000000 992.855000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.140000 0.000000 988.280000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.560000 0.000000 983.700000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.880000 0.000000 979.020000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.305000 0.000000 974.445000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.730000 0.000000 969.870000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.570000 0.000000 965.710000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.995000 0.000000 961.135000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.420000 0.000000 956.560000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.740000 0.000000 951.880000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.160000 0.000000 947.300000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.585000 0.000000 942.725000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.010000 0.000000 938.150000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.330000 0.000000 933.470000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.170000 0.000000 929.310000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.595000 0.000000 924.735000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.120000 0.000000 920.260000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.340000 0.000000 915.480000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.865000 0.000000 911.005000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290000 0.000000 906.430000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.715000 0.000000 901.855000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.140000 0.000000 897.280000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.980000 0.000000 893.120000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.400000 0.000000 888.540000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.825000 0.000000 883.965000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.250000 0.000000 879.390000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.780000 0.000000 874.920000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.995000 0.000000 870.135000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.520000 0.000000 865.660000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.945000 0.000000 861.085000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.785000 0.000000 856.925000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.105000 0.000000 852.245000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.530000 0.000000 847.670000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.955000 0.000000 843.095000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.380000 0.000000 838.520000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.800000 0.000000 833.940000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.120000 0.000000 829.260000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.545000 0.000000 824.685000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.385000 0.000000 820.525000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.810000 0.000000 815.950000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.235000 0.000000 811.375000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.760000 0.000000 806.900000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.980000 0.000000 802.120000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.505000 0.000000 797.645000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.930000 0.000000 793.070000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.355000 0.000000 788.495000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.195000 0.000000 784.335000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.620000 0.000000 779.760000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.040000 0.000000 775.180000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.465000 0.000000 770.605000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.890000 0.000000 766.030000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.210000 0.000000 761.350000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.635000 0.000000 756.775000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.160000 0.000000 752.300000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.000000 0.000000 748.140000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.220000 0.000000 743.360000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.745000 0.000000 738.885000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.170000 0.000000 734.310000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.595000 0.000000 729.735000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.020000 0.000000 725.160000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.340000 0.000000 720.480000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.760000 0.000000 715.900000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.600000 0.000000 711.740000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.025000 0.000000 707.165000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.450000 0.000000 702.590000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.875000 0.000000 698.015000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.195000 0.000000 693.335000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.620000 0.000000 688.760000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.145000 0.000000 684.285000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.570000 0.000000 679.710000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.410000 0.000000 675.550000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.730000 0.000000 670.870000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.155000 0.000000 666.295000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.580000 0.000000 661.720000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.000000 0.000000 657.140000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.320000 0.000000 652.460000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.745000 0.000000 647.885000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170000 0.000000 643.310000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.115000 0.000000 639.255000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.435000 0.000000 634.575000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.860000 0.000000 630.000000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.385000 0.000000 625.525000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.810000 0.000000 620.950000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.235000 0.000000 616.375000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.555000 0.000000 611.695000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.980000 0.000000 607.120000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.920000 0.000000 603.060000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.240000 0.000000 598.380000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.665000 0.000000 593.805000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.090000 0.000000 589.230000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.515000 0.000000 584.655000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.835000 0.000000 579.975000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.260000 0.000000 575.400000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.680000 0.000000 570.820000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.520000 0.000000 566.660000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.840000 0.000000 561.980000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.265000 0.000000 557.405000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.795000 0.000000 552.935000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.148 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2482 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.9455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 548.220000 0.000000 548.360000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0228 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.0535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 543.540000 0.000000 543.680000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.982 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 9.21291 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.804 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 538.960000 0.000000 539.100000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.8212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 534.385000 0.000000 534.525000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.667 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 8.94023 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.9229 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 530.330000 0.000000 530.470000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2998 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.283 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8198 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.8566 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 525.650000 0.000000 525.790000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3053 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 9.28856 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.1707 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 521.075000 0.000000 521.215000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.269 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.6202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 516.500000 0.000000 516.640000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.4405 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8635 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.1484 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 511.920000 0.000000 512.060000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5958 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.2929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 507.450000 0.000000 507.590000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.1545 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 9.58374 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.117 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 502.665000 0.000000 502.805000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4993 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.2805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.737 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.4737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 498.195000 0.000000 498.335000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.402 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 9.50303 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.5222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 493.620000 0.000000 493.760000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.856 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.9204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.2141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 489.460000 0.000000 489.600000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0958 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.37 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 484.780000 0.000000 484.920000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1416 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.364 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.1907 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 480.200000 0.000000 480.340000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1636.370000 0.000000 1636.510000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1631.795000 0.000000 1631.935000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1627.635000 0.000000 1627.775000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1623.060000 0.000000 1623.200000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1618.480000 0.000000 1618.620000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1614.010000 0.000000 1614.150000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1609.435000 0.000000 1609.575000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1604.755000 0.000000 1604.895000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1600.180000 0.000000 1600.320000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1595.600000 0.000000 1595.740000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1591.440000 0.000000 1591.580000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1586.760000 0.000000 1586.900000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1582.185000 0.000000 1582.325000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1577.610000 0.000000 1577.750000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1573.035000 0.000000 1573.175000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1568.355000 0.000000 1568.495000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1563.780000 0.000000 1563.920000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1559.200000 0.000000 1559.340000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1555.040000 0.000000 1555.180000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1550.465000 0.000000 1550.605000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1545.890000 0.000000 1546.030000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1541.210000 0.000000 1541.350000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1536.635000 0.000000 1536.775000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1532.160000 0.000000 1532.300000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1527.585000 0.000000 1527.725000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1523.010000 0.000000 1523.150000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1518.330000 0.000000 1518.470000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1514.275000 0.000000 1514.415000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1509.700000 0.000000 1509.840000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1505.120000 0.000000 1505.260000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1500.545000 0.000000 1500.685000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1495.865000 0.000000 1496.005000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1491.290000 0.000000 1491.430000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1486.820000 0.000000 1486.960000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1482.240000 0.000000 1482.380000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1477.875000 0.000000 1478.015000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1473.400000 0.000000 1473.540000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1468.825000 0.000000 1468.965000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1464.250000 0.000000 1464.390000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1459.675000 0.000000 1459.815000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1454.995000 0.000000 1455.135000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1450.420000 0.000000 1450.560000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1445.840000 0.000000 1445.980000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1441.680000 0.000000 1441.820000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1437.105000 0.000000 1437.245000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1432.425000 0.000000 1432.565000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1427.850000 0.000000 1427.990000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1423.275000 0.000000 1423.415000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1418.800000 0.000000 1418.940000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1414.225000 0.000000 1414.365000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1409.545000 0.000000 1409.685000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1405.385000 0.000000 1405.525000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1400.810000 0.000000 1400.950000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1396.235000 0.000000 1396.375000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1391.555000 0.000000 1391.695000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1386.980000 0.000000 1387.120000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1382.400000 0.000000 1382.540000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1377.825000 0.000000 1377.965000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1373.250000 0.000000 1373.390000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1369.090000 0.000000 1369.230000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1364.515000 0.000000 1364.655000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1360.040000 0.000000 1360.180000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1355.465000 0.000000 1355.605000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1350.890000 0.000000 1351.030000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1346.210000 0.000000 1346.350000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1341.635000 0.000000 1341.775000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1337.060000 0.000000 1337.200000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1332.900000 0.000000 1333.040000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1328.320000 0.000000 1328.460000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1323.640000 0.000000 1323.780000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1319.065000 0.000000 1319.205000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1314.490000 0.000000 1314.630000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1309.915000 0.000000 1310.055000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1305.440000 0.000000 1305.580000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1300.660000 0.000000 1300.800000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1296.500000 0.000000 1296.640000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1292.025000 0.000000 1292.165000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1287.450000 0.000000 1287.590000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1282.770000 0.000000 1282.910000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1278.195000 0.000000 1278.335000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1273.620000 0.000000 1273.760000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1269.040000 0.000000 1269.180000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1264.465000 0.000000 1264.605000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1260.305000 0.000000 1260.445000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1255.730000 0.000000 1255.870000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1251.155000 0.000000 1251.295000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1246.580000 0.000000 1246.720000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1242.105000 0.000000 1242.245000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1237.320000 0.000000 1237.460000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1232.850000 0.000000 1232.990000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1228.275000 0.000000 1228.415000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1224.115000 0.000000 1224.255000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1219.435000 0.000000 1219.575000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1214.860000 0.000000 1215.000000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1210.280000 0.000000 1210.420000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1205.705000 0.000000 1205.845000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1201.130000 0.000000 1201.270000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1196.450000 0.000000 1196.590000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1191.875000 0.000000 1192.015000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1187.715000 0.000000 1187.855000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1183.140000 0.000000 1183.280000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1178.560000 0.000000 1178.700000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1173.880000 0.000000 1174.020000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1169.305000 0.000000 1169.445000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1164.835000 0.000000 1164.975000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1160.260000 0.000000 1160.400000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1155.680000 0.000000 1155.820000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1151.520000 0.000000 1151.660000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1146.945000 0.000000 1147.085000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1142.370000 0.000000 1142.510000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1137.795000 0.000000 1137.935000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1133.220000 0.000000 1133.360000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1128.540000 0.000000 1128.680000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1123.960000 0.000000 1124.100000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1119.490000 0.000000 1119.630000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1115.330000 0.000000 1115.470000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1110.545000 0.000000 1110.685000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1106.075000 0.000000 1106.215000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1101.500000 0.000000 1101.640000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1096.920000 0.000000 1097.060000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1092.345000 0.000000 1092.485000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1087.665000 0.000000 1087.805000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1083.090000 0.000000 1083.230000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1078.930000 0.000000 1079.070000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1074.355000 0.000000 1074.495000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1069.780000 0.000000 1069.920000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1065.100000 0.000000 1065.240000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1060.520000 0.000000 1060.660000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2216.690000 0.000000 2216.830000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.530000 0.000000 2212.670000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2208.060000 0.000000 2208.200000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.480000 0.000000 2203.620000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.800000 0.000000 2198.940000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.225000 0.000000 2194.365000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.650000 0.000000 2189.790000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.075000 0.000000 2185.215000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.395000 0.000000 2180.535000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.340000 0.000000 2176.480000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.760000 0.000000 2171.900000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.080000 0.000000 2167.220000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.505000 0.000000 2162.645000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.930000 0.000000 2158.070000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.460000 0.000000 2153.600000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.880000 0.000000 2149.020000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.200000 0.000000 2144.340000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.040000 0.000000 2140.180000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.465000 0.000000 2135.605000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.890000 0.000000 2131.030000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.210000 0.000000 2126.350000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.635000 0.000000 2121.775000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.060000 0.000000 2117.200000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.480000 0.000000 2112.620000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.905000 0.000000 2108.045000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.745000 0.000000 2103.885000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.170000 0.000000 2099.310000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.700000 0.000000 2094.840000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.120000 0.000000 2090.260000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.440000 0.000000 2085.580000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.865000 0.000000 2081.005000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.290000 0.000000 2076.430000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.610000 0.000000 2071.750000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.555000 0.000000 2067.695000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.980000 0.000000 2063.120000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.300000 0.000000 2058.440000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.720000 0.000000 2053.860000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2049.145000 0.000000 2049.285000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.570000 0.000000 2044.710000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2040.100000 0.000000 2040.240000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.315000 0.000000 2035.455000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.840000 0.000000 2030.980000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.680000 0.000000 2026.820000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.105000 0.000000 2022.245000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.425000 0.000000 2017.565000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.850000 0.000000 2012.990000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.275000 0.000000 2008.415000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.700000 0.000000 2003.840000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.120000 0.000000 1999.260000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.440000 0.000000 1994.580000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.385000 0.000000 1990.525000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.810000 0.000000 1985.950000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.340000 0.000000 1981.480000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.555000 0.000000 1976.695000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.080000 0.000000 1972.220000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.505000 0.000000 1967.645000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.930000 0.000000 1963.070000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.250000 0.000000 1958.390000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.090000 0.000000 1954.230000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.515000 0.000000 1949.655000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.940000 0.000000 1945.080000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.360000 0.000000 1940.500000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.680000 0.000000 1935.820000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.105000 0.000000 1931.245000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.530000 0.000000 1926.670000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.850000 0.000000 1921.990000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.795000 0.000000 1917.935000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.320000 0.000000 1913.460000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.540000 0.000000 1908.680000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.960000 0.000000 1904.100000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.490000 0.000000 1899.630000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.915000 0.000000 1895.055000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.340000 0.000000 1890.480000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.660000 0.000000 1885.800000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.600000 0.000000 1881.740000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.025000 0.000000 1877.165000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.450000 0.000000 1872.590000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.770000 0.000000 1867.910000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.195000 0.000000 1863.335000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.620000 0.000000 1858.760000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.145000 0.000000 1854.285000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.360000 0.000000 1849.500000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.200000 0.000000 1845.340000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.730000 0.000000 1840.870000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.155000 0.000000 1836.295000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.580000 0.000000 1831.720000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.900000 0.000000 1827.040000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.320000 0.000000 1822.460000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.745000 0.000000 1817.885000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.170000 0.000000 1813.310000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.010000 0.000000 1809.150000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.435000 0.000000 1804.575000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.755000 0.000000 1799.895000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.180000 0.000000 1795.320000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.600000 0.000000 1790.740000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.130000 0.000000 1786.270000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.555000 0.000000 1781.695000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.875000 0.000000 1777.015000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.715000 0.000000 1772.855000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.140000 0.000000 1768.280000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.560000 0.000000 1763.700000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.880000 0.000000 1759.020000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.305000 0.000000 1754.445000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.730000 0.000000 1749.870000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.155000 0.000000 1745.295000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.580000 0.000000 1740.720000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.420000 0.000000 1736.560000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.840000 0.000000 1731.980000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.370000 0.000000 1727.510000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.795000 0.000000 1722.935000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.115000 0.000000 1718.255000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.540000 0.000000 1713.680000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.960000 0.000000 1709.100000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.385000 0.000000 1704.525000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.225000 0.000000 1700.365000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.650000 0.000000 1695.790000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.970000 0.000000 1691.110000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.395000 0.000000 1686.535000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.820000 0.000000 1681.960000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.240000 0.000000 1677.380000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.770000 0.000000 1672.910000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.985000 0.000000 1668.125000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.825000 0.000000 1663.965000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1659.355000 0.000000 1659.495000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.780000 0.000000 1654.920000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.100000 0.000000 1650.240000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.520000 0.000000 1645.660000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.945000 0.000000 1641.085000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 77.450000 0.800000 77.750000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 183.913 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 982.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.731 LAYER met4  ;
    ANTENNAMAXAREACAR 161.169 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 854.919 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.394653 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.050000 0.800000 194.350000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 166.648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 890.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.731 LAYER met4  ;
    ANTENNAMAXAREACAR 146.031 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 761.582 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.340013 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 310.950000 0.800000 311.250000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 116.895 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 625.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4705 LAYER met4  ;
    ANTENNAMAXAREACAR 65.6972 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 345.282 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.385484 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 466.150000 0.800000 466.450000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.4944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 312.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 65.6226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 353.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 55.8301 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.939 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 621.550000 0.800000 621.850000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 776.950000 0.800000 777.250000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 932.750000 0.800000 933.050000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1088.250000 0.800000 1088.550000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 29.5401 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 155.183 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 0.5644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.472 LAYER met3  ;
    ANTENNAGATEAREA 0.9366 LAYER met3  ;
    ANTENNAMAXAREACAR 77.4279 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 369.599 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.629216 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1243.550000 0.800000 1243.850000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 26.5218 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 139.981 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 2.1193 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.768 LAYER met3  ;
    ANTENNAGATEAREA 0.9366 LAYER met3  ;
    ANTENNAMAXAREACAR 49.8986 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 233.368 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.450644 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1398.750000 0.800000 1399.050000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 43.4833 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 196.762 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1554.650000 0.800000 1554.950000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 64.6613 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 322.671 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1710.050000 0.800000 1710.350000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 39.6302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 197.135 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 61.8454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 330.304 LAYER met3  ;
    ANTENNAGATEAREA 0.9366 LAYER met3  ;
    ANTENNAMAXAREACAR 140.88 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 724.249 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.450644 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1865.450000 0.800000 1865.750000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9742 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 17.2561 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.8779 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2020.950000 0.800000 2021.250000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.1795 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 60.1506 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 297.313 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 127.640000 2118.390000 127.780000 2118.880000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.0875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 60.3829 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 299.62 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 383.275000 2118.390000 383.415000 2118.880000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 101.721 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 522.865 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 46.5178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 232.428 LAYER met2  ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 90.026 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 422.361 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 638.595000 2118.390000 638.735000 2118.880000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 45.8357 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.786 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 12.7526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.602 LAYER met2  ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 75.8347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 362.42 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.480404 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 894.435000 2118.390000 894.575000 2118.880000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.0475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 42.5049 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 210.23 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1149.650000 2118.390000 1149.790000 2118.880000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.6955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 36.9384 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 181.252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1404.970000 2118.390000 1405.110000 2118.880000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7437 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 250.452 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 32.0005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 159.842 LAYER met2  ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 79.2167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 369.355 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.396032 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1660.810000 2118.390000 1660.950000 2118.880000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 102.914 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 529.365 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 6.0681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0615 LAYER met2  ;
    ANTENNAGATEAREA 0.9366 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4196 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 318.909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1915.920000 2118.390000 1916.060000 2118.880000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 64.8135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 308.845 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.6584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.066 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 34.7737 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.641 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.580051 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2171.760000 2118.390000 2171.900000 2118.880000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 80.0601 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 397.653 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1979.950000 2299.540000 1980.250000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 168.306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 898.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 62.0413 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 324.794 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1821.750000 2299.540000 1822.050000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 121.257 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 647.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 76.3842 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 415.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1663.350000 2299.540000 1663.650000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.3306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.1554 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 108.358 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 542.615 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1504.650000 2299.540000 1504.950000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6013 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met4  ;
    ANTENNAMAXAREACAR 27.7134 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.653 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616901 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1346.250000 2299.540000 1346.550000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1187.850000 2299.540000 1188.150000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1029.550000 2299.540000 1029.850000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 575.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.95 LAYER met3  ;
    ANTENNAMAXAREACAR 82.6356 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 415.751 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.408509 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 870.750000 2299.540000 871.050000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 712.450000 2299.540000 712.750000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 127.292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 678.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.72 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.192 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285 LAYER met4  ;
    ANTENNAMAXAREACAR 75.6931 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.462 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 593.550000 2299.540000 593.850000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 474.750000 2299.540000 475.050000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 355.750000 2299.540000 356.050000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 151.245 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 807.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.5758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 71.025 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 374.865 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 236.950000 2299.540000 237.250000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 118.050000 2299.540000 118.350000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 2.750000 2299.540000 3.050000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 839.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 38.750000 0.800000 39.050000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.550000 0.800000 155.850000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 271.750000 0.800000 272.050000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.1534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 427.250000 0.800000 427.550000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 583.050000 0.800000 583.350000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 738.450000 0.800000 738.750000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 300.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1604.93 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 112.594 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 601.44 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 893.750000 0.800000 894.050000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.276 LAYER met3  ;
    ANTENNAMAXAREACAR 80.6557 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 399.992 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.280067 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1049.050000 0.800000 1049.350000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.801 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 33.6158 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.081 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1204.850000 0.800000 1205.150000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 70.8848 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 378.952 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854141 LAYER via4  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.176 LAYER met3  ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 61.6175 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 323.203 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1360.350000 0.800000 1360.650000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.4164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 5.1422 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.674 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 166.111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 904.57 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854141 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1515.750000 0.800000 1516.050000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1670.950000 0.800000 1671.250000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1826.450000 0.800000 1826.750000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1982.150000 0.800000 1982.450000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.5265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.785000 2118.390000 63.925000 2118.880000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 65.8018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 328.783 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 319.420000 2118.390000 319.560000 2118.880000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 60.5392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 302.47 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 574.840000 2118.390000 574.980000 2118.880000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.5613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 292.646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.1868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 49.4327 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 256.504 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.261549 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 830.060000 2118.390000 830.200000 2118.880000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 59.3506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 296.527 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1085.900000 2118.390000 1086.040000 2118.880000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 63.9768 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 319.648 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 259.935 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 1297.13 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1341.115000 2118.390000 1341.255000 2118.880000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 58.2019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 290.783 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1596.955000 2118.390000 1597.095000 2118.880000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 66.2933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 330.887 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 92.7819 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 461.107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1852.065000 2118.390000 1852.205000 2118.880000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 29.9848 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.383 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 59.9219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 299.331 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.16 LAYER met3  ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 28.5925 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 139.324 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.404646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2107.905000 2118.390000 2108.045000 2118.880000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.36 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 2019.550000 2299.540000 2019.850000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.8976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.728 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1861.250000 2299.540000 1861.550000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 372.911 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1989.79 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1702.850000 2299.540000 1703.150000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 40.2522 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 215.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1544.550000 2299.540000 1544.850000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.7102 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1385.650000 2299.540000 1385.950000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1227.350000 2299.540000 1227.650000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1069.050000 2299.540000 1069.350000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.375 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 910.650000 2299.540000 910.950000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 253.545 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1353.18 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 751.950000 2299.540000 752.250000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.375 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 633.050000 2299.540000 633.350000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 514.250000 2299.540000 514.550000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.3834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 395.750000 2299.540000 396.050000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 839.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 276.950000 2299.540000 277.250000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 158.050000 2299.540000 158.350000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 96.3184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 514.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.5808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 339.568 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 39.250000 2299.540000 39.550000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 839.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 3.550000 0.800000 3.850000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.0254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.450000 0.800000 116.750000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 233.250000 0.800000 233.550000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 388.550000 0.800000 388.850000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 543.950000 0.800000 544.250000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 839.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 699.250000 0.800000 699.550000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 839.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 855.050000 0.800000 855.350000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 839.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1010.550000 0.800000 1010.850000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1165.750000 0.800000 1166.050000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.2862 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.992 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1321.250000 0.800000 1321.550000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.4722 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.984 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1476.550000 0.800000 1476.850000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1632.350000 0.800000 1632.650000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 41.4252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 221.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1787.850000 0.800000 1788.150000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1943.150000 0.800000 1943.450000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.0679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.2115 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.025000 2118.390000 5.165000 2118.880000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.0778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 320.11 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.08 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 255.145000 2118.390000 255.285000 2118.880000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 57.0791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 285.169 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 510.985000 2118.390000 511.125000 2118.880000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 53.8514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 269.031 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 766.200000 2118.390000 766.340000 2118.880000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 59.2421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 295.984 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1022.040000 2118.390000 1022.180000 2118.880000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 57.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 288.295 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1277.260000 2118.390000 1277.400000 2118.880000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 58.4406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 291.977 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1533.100000 2118.390000 1533.240000 2118.880000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6626 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 53.5238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 267.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1788.420000 2118.390000 1788.560000 2118.880000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 64.2918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 320.761 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2044.050000 2118.390000 2044.190000 2118.880000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 2055.650000 2299.540000 2055.950000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 240.283 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1281.98 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1901.050000 2299.540000 1901.350000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1742.350000 2299.540000 1742.650000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1584.050000 2299.540000 1584.350000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1425.650000 2299.540000 1425.950000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.4574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1266.850000 2299.540000 1267.150000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1108.550000 2299.540000 1108.850000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4982 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 950.050000 2299.540000 950.350000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.375 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 791.850000 2299.540000 792.150000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4982 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 672.950000 2299.540000 673.250000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.375 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 554.150000 2299.540000 554.450000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.375 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 435.150000 2299.540000 435.450000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4532 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 316.450000 2299.540000 316.750000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.3854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.384 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 197.450000 2299.540000 197.750000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.375 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 78.650000 2299.540000 78.950000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 349.450000 0.800000 349.750000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 505.350000 0.800000 505.650000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 660.750000 0.800000 661.050000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 816.050000 0.800000 816.350000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 971.250000 0.800000 971.550000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1126.750000 0.800000 1127.050000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1282.550000 0.800000 1282.850000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1437.950000 0.800000 1438.250000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1593.450000 0.800000 1593.750000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1748.750000 0.800000 1749.050000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1904.450000 0.800000 1904.750000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2056.350000 0.800000 2056.650000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.500000 2118.390000 191.640000 2118.880000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.130000 2118.390000 447.270000 2118.880000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.450000 2118.390000 702.590000 2118.880000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.185000 2118.390000 958.325000 2118.880000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.610000 2118.390000 1213.750000 2118.880000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.240000 2118.390000 1469.380000 2118.880000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.460000 2118.390000 1724.600000 2118.880000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.780000 2118.390000 1979.920000 2118.880000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.940000 2118.390000 2231.080000 2118.880000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1940.550000 2299.540000 1940.850000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1782.150000 2299.540000 1782.450000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1623.450000 2299.540000 1623.750000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1465.050000 2299.540000 1465.350000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1306.750000 2299.540000 1307.050000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 1148.450000 2299.540000 1148.750000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 989.750000 2299.540000 990.050000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2298.740000 831.350000 2299.540000 831.650000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.265000 0.000000 2221.405000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.669 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2235.100000 0.000000 2235.240000 0.490000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.77 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2230.520000 0.000000 2230.660000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.522 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 156.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 840.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2225.945000 0.000000 2226.085000 0.490000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2276.520000 13.120000 2286.520000 2104.400000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.020000 13.120000 23.020000 2104.400000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 538.400000 170.660000 540.140000 565.440000 ;
      LAYER met3 ;
        RECT 63.080000 170.660000 540.140000 172.400000 ;
      LAYER met3 ;
        RECT 63.080000 563.700000 540.140000 565.440000 ;
      LAYER met4 ;
        RECT 63.080000 170.660000 64.820000 565.440000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 538.400000 668.160000 540.140000 1062.940000 ;
      LAYER met3 ;
        RECT 63.080000 668.160000 540.140000 669.900000 ;
      LAYER met3 ;
        RECT 63.080000 1061.200000 540.140000 1062.940000 ;
      LAYER met4 ;
        RECT 63.080000 668.160000 64.820000 1062.940000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 538.400000 1165.660000 540.140000 1560.440000 ;
      LAYER met3 ;
        RECT 63.080000 1165.660000 540.140000 1167.400000 ;
      LAYER met3 ;
        RECT 63.080000 1558.700000 540.140000 1560.440000 ;
      LAYER met4 ;
        RECT 63.080000 1165.660000 64.820000 1560.440000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 538.400000 1663.160000 540.140000 2057.940000 ;
      LAYER met3 ;
        RECT 63.080000 1663.160000 540.140000 1664.900000 ;
      LAYER met3 ;
        RECT 63.080000 2056.200000 540.140000 2057.940000 ;
      LAYER met4 ;
        RECT 63.080000 1663.160000 64.820000 2057.940000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2238.180000 170.660000 2239.920000 565.440000 ;
      LAYER met3 ;
        RECT 1762.860000 170.660000 2239.920000 172.400000 ;
      LAYER met3 ;
        RECT 1762.860000 563.700000 2239.920000 565.440000 ;
      LAYER met4 ;
        RECT 1762.860000 170.660000 1764.600000 565.440000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2238.180000 668.160000 2239.920000 1062.940000 ;
      LAYER met3 ;
        RECT 1762.860000 668.160000 2239.920000 669.900000 ;
      LAYER met3 ;
        RECT 1762.860000 1061.200000 2239.920000 1062.940000 ;
      LAYER met4 ;
        RECT 1762.860000 668.160000 1764.600000 1062.940000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2238.180000 1165.660000 2239.920000 1560.440000 ;
      LAYER met3 ;
        RECT 1762.860000 1165.660000 2239.920000 1167.400000 ;
      LAYER met3 ;
        RECT 1762.860000 1558.700000 2239.920000 1560.440000 ;
      LAYER met4 ;
        RECT 1762.860000 1165.660000 1764.600000 1560.440000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2238.180000 1663.160000 2239.920000 2057.940000 ;
      LAYER met3 ;
        RECT 1762.860000 1663.160000 2239.920000 1664.900000 ;
      LAYER met3 ;
        RECT 1762.860000 2056.200000 2239.920000 2057.940000 ;
      LAYER met4 ;
        RECT 1762.860000 1663.160000 1764.600000 2057.940000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2264.520000 25.120000 2274.520000 2092.400000 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.020000 25.120000 35.020000 2092.400000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 66.480000 560.300000 536.740000 562.040000 ;
      LAYER met3 ;
        RECT 66.480000 174.060000 536.740000 175.800000 ;
      LAYER met4 ;
        RECT 66.480000 174.060000 68.220000 562.040000 ;
      LAYER met4 ;
        RECT 535.000000 174.060000 536.740000 562.040000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 66.480000 1057.800000 536.740000 1059.540000 ;
      LAYER met3 ;
        RECT 66.480000 671.560000 536.740000 673.300000 ;
      LAYER met4 ;
        RECT 66.480000 671.560000 68.220000 1059.540000 ;
      LAYER met4 ;
        RECT 535.000000 671.560000 536.740000 1059.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 66.480000 1555.300000 536.740000 1557.040000 ;
      LAYER met3 ;
        RECT 66.480000 1169.060000 536.740000 1170.800000 ;
      LAYER met4 ;
        RECT 66.480000 1169.060000 68.220000 1557.040000 ;
      LAYER met4 ;
        RECT 535.000000 1169.060000 536.740000 1557.040000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 66.480000 2052.800000 536.740000 2054.540000 ;
      LAYER met3 ;
        RECT 66.480000 1666.560000 536.740000 1668.300000 ;
      LAYER met4 ;
        RECT 66.480000 1666.560000 68.220000 2054.540000 ;
      LAYER met4 ;
        RECT 535.000000 1666.560000 536.740000 2054.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1766.260000 560.300000 2236.520000 562.040000 ;
      LAYER met3 ;
        RECT 1766.260000 174.060000 2236.520000 175.800000 ;
      LAYER met4 ;
        RECT 1766.260000 174.060000 1768.000000 562.040000 ;
      LAYER met4 ;
        RECT 2234.780000 174.060000 2236.520000 562.040000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1766.260000 1057.800000 2236.520000 1059.540000 ;
      LAYER met3 ;
        RECT 1766.260000 671.560000 2236.520000 673.300000 ;
      LAYER met4 ;
        RECT 1766.260000 671.560000 1768.000000 1059.540000 ;
      LAYER met4 ;
        RECT 2234.780000 671.560000 2236.520000 1059.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1766.260000 1555.300000 2236.520000 1557.040000 ;
      LAYER met3 ;
        RECT 1766.260000 1169.060000 2236.520000 1170.800000 ;
      LAYER met4 ;
        RECT 1766.260000 1169.060000 1768.000000 1557.040000 ;
      LAYER met4 ;
        RECT 2234.780000 1169.060000 2236.520000 1557.040000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1766.260000 2052.800000 2236.520000 2054.540000 ;
      LAYER met3 ;
        RECT 1766.260000 1666.560000 2236.520000 1668.300000 ;
      LAYER met4 ;
        RECT 1766.260000 1666.560000 1768.000000 2054.540000 ;
      LAYER met4 ;
        RECT 2234.780000 1666.560000 2236.520000 2054.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2299.540000 2118.880000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2299.540000 2118.880000 ;
    LAYER met2 ;
      RECT 2231.220000 2118.250000 2299.540000 2118.880000 ;
      RECT 2172.040000 2118.250000 2230.800000 2118.880000 ;
      RECT 2108.185000 2118.250000 2171.620000 2118.880000 ;
      RECT 2044.330000 2118.250000 2107.765000 2118.880000 ;
      RECT 1980.060000 2118.250000 2043.910000 2118.880000 ;
      RECT 1916.200000 2118.250000 1979.640000 2118.880000 ;
      RECT 1852.345000 2118.250000 1915.780000 2118.880000 ;
      RECT 1788.700000 2118.250000 1851.925000 2118.880000 ;
      RECT 1724.740000 2118.250000 1788.280000 2118.880000 ;
      RECT 1661.090000 2118.250000 1724.320000 2118.880000 ;
      RECT 1597.235000 2118.250000 1660.670000 2118.880000 ;
      RECT 1533.380000 2118.250000 1596.815000 2118.880000 ;
      RECT 1469.520000 2118.250000 1532.960000 2118.880000 ;
      RECT 1405.250000 2118.250000 1469.100000 2118.880000 ;
      RECT 1341.395000 2118.250000 1404.830000 2118.880000 ;
      RECT 1277.540000 2118.250000 1340.975000 2118.880000 ;
      RECT 1213.890000 2118.250000 1277.120000 2118.880000 ;
      RECT 1149.930000 2118.250000 1213.470000 2118.880000 ;
      RECT 1086.180000 2118.250000 1149.510000 2118.880000 ;
      RECT 1022.320000 2118.250000 1085.760000 2118.880000 ;
      RECT 958.465000 2118.250000 1021.900000 2118.880000 ;
      RECT 894.715000 2118.250000 958.045000 2118.880000 ;
      RECT 830.340000 2118.250000 894.295000 2118.880000 ;
      RECT 766.480000 2118.250000 829.920000 2118.880000 ;
      RECT 702.730000 2118.250000 766.060000 2118.880000 ;
      RECT 638.875000 2118.250000 702.310000 2118.880000 ;
      RECT 575.120000 2118.250000 638.455000 2118.880000 ;
      RECT 511.265000 2118.250000 574.700000 2118.880000 ;
      RECT 447.410000 2118.250000 510.845000 2118.880000 ;
      RECT 383.555000 2118.250000 446.990000 2118.880000 ;
      RECT 319.700000 2118.250000 383.135000 2118.880000 ;
      RECT 255.425000 2118.250000 319.280000 2118.880000 ;
      RECT 191.780000 2118.250000 255.005000 2118.880000 ;
      RECT 127.920000 2118.250000 191.360000 2118.880000 ;
      RECT 64.065000 2118.250000 127.500000 2118.880000 ;
      RECT 5.305000 2118.250000 63.645000 2118.880000 ;
      RECT 0.000000 2118.250000 4.885000 2118.880000 ;
      RECT 0.000000 0.630000 2299.540000 2118.250000 ;
      RECT 4.370000 0.625000 8.420000 0.630000 ;
      RECT 2235.380000 0.000000 2299.540000 0.630000 ;
      RECT 2230.800000 0.000000 2234.960000 0.630000 ;
      RECT 2226.225000 0.000000 2230.380000 0.630000 ;
      RECT 2221.545000 0.000000 2225.805000 0.630000 ;
      RECT 2216.970000 0.000000 2221.125000 0.630000 ;
      RECT 2212.810000 0.000000 2216.550000 0.630000 ;
      RECT 2208.340000 0.000000 2212.390000 0.630000 ;
      RECT 2203.760000 0.000000 2207.920000 0.630000 ;
      RECT 2199.080000 0.000000 2203.340000 0.630000 ;
      RECT 2194.505000 0.000000 2198.660000 0.630000 ;
      RECT 2189.930000 0.000000 2194.085000 0.630000 ;
      RECT 2185.355000 0.000000 2189.510000 0.630000 ;
      RECT 2180.675000 0.000000 2184.935000 0.630000 ;
      RECT 2176.620000 0.000000 2180.255000 0.630000 ;
      RECT 2172.040000 0.000000 2176.200000 0.630000 ;
      RECT 2167.360000 0.000000 2171.620000 0.630000 ;
      RECT 2162.785000 0.000000 2166.940000 0.630000 ;
      RECT 2158.210000 0.000000 2162.365000 0.630000 ;
      RECT 2153.740000 0.000000 2157.790000 0.630000 ;
      RECT 2149.160000 0.000000 2153.320000 0.630000 ;
      RECT 2144.480000 0.000000 2148.740000 0.630000 ;
      RECT 2140.320000 0.000000 2144.060000 0.630000 ;
      RECT 2135.745000 0.000000 2139.900000 0.630000 ;
      RECT 2131.170000 0.000000 2135.325000 0.630000 ;
      RECT 2126.490000 0.000000 2130.750000 0.630000 ;
      RECT 2121.915000 0.000000 2126.070000 0.630000 ;
      RECT 2117.340000 0.000000 2121.495000 0.630000 ;
      RECT 2112.760000 0.000000 2116.920000 0.630000 ;
      RECT 2108.185000 0.000000 2112.340000 0.630000 ;
      RECT 2104.025000 0.000000 2107.765000 0.630000 ;
      RECT 2099.450000 0.000000 2103.605000 0.630000 ;
      RECT 2094.980000 0.000000 2099.030000 0.630000 ;
      RECT 2090.400000 0.000000 2094.560000 0.630000 ;
      RECT 2085.720000 0.000000 2089.980000 0.630000 ;
      RECT 2081.145000 0.000000 2085.300000 0.630000 ;
      RECT 2076.570000 0.000000 2080.725000 0.630000 ;
      RECT 2071.890000 0.000000 2076.150000 0.630000 ;
      RECT 2067.835000 0.000000 2071.470000 0.630000 ;
      RECT 2063.260000 0.000000 2067.415000 0.630000 ;
      RECT 2058.580000 0.000000 2062.840000 0.630000 ;
      RECT 2054.000000 0.000000 2058.160000 0.630000 ;
      RECT 2049.425000 0.000000 2053.580000 0.630000 ;
      RECT 2044.850000 0.000000 2049.005000 0.630000 ;
      RECT 2040.380000 0.000000 2044.430000 0.630000 ;
      RECT 2035.595000 0.000000 2039.960000 0.630000 ;
      RECT 2031.120000 0.000000 2035.175000 0.630000 ;
      RECT 2026.960000 0.000000 2030.700000 0.630000 ;
      RECT 2022.385000 0.000000 2026.540000 0.630000 ;
      RECT 2017.705000 0.000000 2021.965000 0.630000 ;
      RECT 2013.130000 0.000000 2017.285000 0.630000 ;
      RECT 2008.555000 0.000000 2012.710000 0.630000 ;
      RECT 2003.980000 0.000000 2008.135000 0.630000 ;
      RECT 1999.400000 0.000000 2003.560000 0.630000 ;
      RECT 1994.720000 0.000000 1998.980000 0.630000 ;
      RECT 1990.665000 0.000000 1994.300000 0.630000 ;
      RECT 1986.090000 0.000000 1990.245000 0.630000 ;
      RECT 1981.620000 0.000000 1985.670000 0.630000 ;
      RECT 1976.835000 0.000000 1981.200000 0.630000 ;
      RECT 1972.360000 0.000000 1976.415000 0.630000 ;
      RECT 1967.785000 0.000000 1971.940000 0.630000 ;
      RECT 1963.210000 0.000000 1967.365000 0.630000 ;
      RECT 1958.530000 0.000000 1962.790000 0.630000 ;
      RECT 1954.370000 0.000000 1958.110000 0.630000 ;
      RECT 1949.795000 0.000000 1953.950000 0.630000 ;
      RECT 1945.220000 0.000000 1949.375000 0.630000 ;
      RECT 1940.640000 0.000000 1944.800000 0.630000 ;
      RECT 1935.960000 0.000000 1940.220000 0.630000 ;
      RECT 1931.385000 0.000000 1935.540000 0.630000 ;
      RECT 1926.810000 0.000000 1930.965000 0.630000 ;
      RECT 1922.130000 0.000000 1926.390000 0.630000 ;
      RECT 1918.075000 0.000000 1921.710000 0.630000 ;
      RECT 1913.600000 0.000000 1917.655000 0.630000 ;
      RECT 1908.820000 0.000000 1913.180000 0.630000 ;
      RECT 1904.240000 0.000000 1908.400000 0.630000 ;
      RECT 1899.770000 0.000000 1903.820000 0.630000 ;
      RECT 1895.195000 0.000000 1899.350000 0.630000 ;
      RECT 1890.620000 0.000000 1894.775000 0.630000 ;
      RECT 1885.940000 0.000000 1890.200000 0.630000 ;
      RECT 1881.880000 0.000000 1885.520000 0.630000 ;
      RECT 1877.305000 0.000000 1881.460000 0.630000 ;
      RECT 1872.730000 0.000000 1876.885000 0.630000 ;
      RECT 1868.050000 0.000000 1872.310000 0.630000 ;
      RECT 1863.475000 0.000000 1867.630000 0.630000 ;
      RECT 1858.900000 0.000000 1863.055000 0.630000 ;
      RECT 1854.425000 0.000000 1858.480000 0.630000 ;
      RECT 1849.640000 0.000000 1854.005000 0.630000 ;
      RECT 1845.480000 0.000000 1849.220000 0.630000 ;
      RECT 1841.010000 0.000000 1845.060000 0.630000 ;
      RECT 1836.435000 0.000000 1840.590000 0.630000 ;
      RECT 1831.860000 0.000000 1836.015000 0.630000 ;
      RECT 1827.180000 0.000000 1831.440000 0.630000 ;
      RECT 1822.600000 0.000000 1826.760000 0.630000 ;
      RECT 1818.025000 0.000000 1822.180000 0.630000 ;
      RECT 1813.450000 0.000000 1817.605000 0.630000 ;
      RECT 1809.290000 0.000000 1813.030000 0.630000 ;
      RECT 1804.715000 0.000000 1808.870000 0.630000 ;
      RECT 1800.035000 0.000000 1804.295000 0.630000 ;
      RECT 1795.460000 0.000000 1799.615000 0.630000 ;
      RECT 1790.880000 0.000000 1795.040000 0.630000 ;
      RECT 1786.410000 0.000000 1790.460000 0.630000 ;
      RECT 1781.835000 0.000000 1785.990000 0.630000 ;
      RECT 1777.155000 0.000000 1781.415000 0.630000 ;
      RECT 1772.995000 0.000000 1776.735000 0.630000 ;
      RECT 1768.420000 0.000000 1772.575000 0.630000 ;
      RECT 1763.840000 0.000000 1768.000000 0.630000 ;
      RECT 1759.160000 0.000000 1763.420000 0.630000 ;
      RECT 1754.585000 0.000000 1758.740000 0.630000 ;
      RECT 1750.010000 0.000000 1754.165000 0.630000 ;
      RECT 1745.435000 0.000000 1749.590000 0.630000 ;
      RECT 1740.860000 0.000000 1745.015000 0.630000 ;
      RECT 1736.700000 0.000000 1740.440000 0.630000 ;
      RECT 1732.120000 0.000000 1736.280000 0.630000 ;
      RECT 1727.650000 0.000000 1731.700000 0.630000 ;
      RECT 1723.075000 0.000000 1727.230000 0.630000 ;
      RECT 1718.395000 0.000000 1722.655000 0.630000 ;
      RECT 1713.820000 0.000000 1717.975000 0.630000 ;
      RECT 1709.240000 0.000000 1713.400000 0.630000 ;
      RECT 1704.665000 0.000000 1708.820000 0.630000 ;
      RECT 1700.505000 0.000000 1704.245000 0.630000 ;
      RECT 1695.930000 0.000000 1700.085000 0.630000 ;
      RECT 1691.250000 0.000000 1695.510000 0.630000 ;
      RECT 1686.675000 0.000000 1690.830000 0.630000 ;
      RECT 1682.100000 0.000000 1686.255000 0.630000 ;
      RECT 1677.520000 0.000000 1681.680000 0.630000 ;
      RECT 1673.050000 0.000000 1677.100000 0.630000 ;
      RECT 1668.265000 0.000000 1672.630000 0.630000 ;
      RECT 1664.105000 0.000000 1667.845000 0.630000 ;
      RECT 1659.635000 0.000000 1663.685000 0.630000 ;
      RECT 1655.060000 0.000000 1659.215000 0.630000 ;
      RECT 1650.380000 0.000000 1654.640000 0.630000 ;
      RECT 1645.800000 0.000000 1649.960000 0.630000 ;
      RECT 1641.225000 0.000000 1645.380000 0.630000 ;
      RECT 1636.650000 0.000000 1640.805000 0.630000 ;
      RECT 1632.075000 0.000000 1636.230000 0.630000 ;
      RECT 1627.915000 0.000000 1631.655000 0.630000 ;
      RECT 1623.340000 0.000000 1627.495000 0.630000 ;
      RECT 1618.760000 0.000000 1622.920000 0.630000 ;
      RECT 1614.290000 0.000000 1618.340000 0.630000 ;
      RECT 1609.715000 0.000000 1613.870000 0.630000 ;
      RECT 1605.035000 0.000000 1609.295000 0.630000 ;
      RECT 1600.460000 0.000000 1604.615000 0.630000 ;
      RECT 1595.880000 0.000000 1600.040000 0.630000 ;
      RECT 1591.720000 0.000000 1595.460000 0.630000 ;
      RECT 1587.040000 0.000000 1591.300000 0.630000 ;
      RECT 1582.465000 0.000000 1586.620000 0.630000 ;
      RECT 1577.890000 0.000000 1582.045000 0.630000 ;
      RECT 1573.315000 0.000000 1577.470000 0.630000 ;
      RECT 1568.635000 0.000000 1572.895000 0.630000 ;
      RECT 1564.060000 0.000000 1568.215000 0.630000 ;
      RECT 1559.480000 0.000000 1563.640000 0.630000 ;
      RECT 1555.320000 0.000000 1559.060000 0.630000 ;
      RECT 1550.745000 0.000000 1554.900000 0.630000 ;
      RECT 1546.170000 0.000000 1550.325000 0.630000 ;
      RECT 1541.490000 0.000000 1545.750000 0.630000 ;
      RECT 1536.915000 0.000000 1541.070000 0.630000 ;
      RECT 1532.440000 0.000000 1536.495000 0.630000 ;
      RECT 1527.865000 0.000000 1532.020000 0.630000 ;
      RECT 1523.290000 0.000000 1527.445000 0.630000 ;
      RECT 1518.610000 0.000000 1522.870000 0.630000 ;
      RECT 1514.555000 0.000000 1518.190000 0.630000 ;
      RECT 1509.980000 0.000000 1514.135000 0.630000 ;
      RECT 1505.400000 0.000000 1509.560000 0.630000 ;
      RECT 1500.825000 0.000000 1504.980000 0.630000 ;
      RECT 1496.145000 0.000000 1500.405000 0.630000 ;
      RECT 1491.570000 0.000000 1495.725000 0.630000 ;
      RECT 1487.100000 0.000000 1491.150000 0.630000 ;
      RECT 1482.520000 0.000000 1486.680000 0.630000 ;
      RECT 1478.155000 0.000000 1482.100000 0.630000 ;
      RECT 1473.680000 0.000000 1477.735000 0.630000 ;
      RECT 1469.105000 0.000000 1473.260000 0.630000 ;
      RECT 1464.530000 0.000000 1468.685000 0.630000 ;
      RECT 1459.955000 0.000000 1464.110000 0.630000 ;
      RECT 1455.275000 0.000000 1459.535000 0.630000 ;
      RECT 1450.700000 0.000000 1454.855000 0.630000 ;
      RECT 1446.120000 0.000000 1450.280000 0.630000 ;
      RECT 1441.960000 0.000000 1445.700000 0.630000 ;
      RECT 1437.385000 0.000000 1441.540000 0.630000 ;
      RECT 1432.705000 0.000000 1436.965000 0.630000 ;
      RECT 1428.130000 0.000000 1432.285000 0.630000 ;
      RECT 1423.555000 0.000000 1427.710000 0.630000 ;
      RECT 1419.080000 0.000000 1423.135000 0.630000 ;
      RECT 1414.505000 0.000000 1418.660000 0.630000 ;
      RECT 1409.825000 0.000000 1414.085000 0.630000 ;
      RECT 1405.665000 0.000000 1409.405000 0.630000 ;
      RECT 1401.090000 0.000000 1405.245000 0.630000 ;
      RECT 1396.515000 0.000000 1400.670000 0.630000 ;
      RECT 1391.835000 0.000000 1396.095000 0.630000 ;
      RECT 1387.260000 0.000000 1391.415000 0.630000 ;
      RECT 1382.680000 0.000000 1386.840000 0.630000 ;
      RECT 1378.105000 0.000000 1382.260000 0.630000 ;
      RECT 1373.530000 0.000000 1377.685000 0.630000 ;
      RECT 1369.370000 0.000000 1373.110000 0.630000 ;
      RECT 1364.795000 0.000000 1368.950000 0.630000 ;
      RECT 1360.320000 0.000000 1364.375000 0.630000 ;
      RECT 1355.745000 0.000000 1359.900000 0.630000 ;
      RECT 1351.170000 0.000000 1355.325000 0.630000 ;
      RECT 1346.490000 0.000000 1350.750000 0.630000 ;
      RECT 1341.915000 0.000000 1346.070000 0.630000 ;
      RECT 1337.340000 0.000000 1341.495000 0.630000 ;
      RECT 1333.180000 0.000000 1336.920000 0.630000 ;
      RECT 1328.600000 0.000000 1332.760000 0.630000 ;
      RECT 1323.920000 0.000000 1328.180000 0.630000 ;
      RECT 1319.345000 0.000000 1323.500000 0.630000 ;
      RECT 1314.770000 0.000000 1318.925000 0.630000 ;
      RECT 1310.195000 0.000000 1314.350000 0.630000 ;
      RECT 1305.720000 0.000000 1309.775000 0.630000 ;
      RECT 1300.940000 0.000000 1305.300000 0.630000 ;
      RECT 1296.780000 0.000000 1300.520000 0.630000 ;
      RECT 1292.305000 0.000000 1296.360000 0.630000 ;
      RECT 1287.730000 0.000000 1291.885000 0.630000 ;
      RECT 1283.050000 0.000000 1287.310000 0.630000 ;
      RECT 1278.475000 0.000000 1282.630000 0.630000 ;
      RECT 1273.900000 0.000000 1278.055000 0.630000 ;
      RECT 1269.320000 0.000000 1273.480000 0.630000 ;
      RECT 1264.745000 0.000000 1268.900000 0.630000 ;
      RECT 1260.585000 0.000000 1264.325000 0.630000 ;
      RECT 1256.010000 0.000000 1260.165000 0.630000 ;
      RECT 1251.435000 0.000000 1255.590000 0.630000 ;
      RECT 1246.860000 0.000000 1251.015000 0.630000 ;
      RECT 1242.385000 0.000000 1246.440000 0.630000 ;
      RECT 1237.600000 0.000000 1241.965000 0.630000 ;
      RECT 1233.130000 0.000000 1237.180000 0.630000 ;
      RECT 1228.555000 0.000000 1232.710000 0.630000 ;
      RECT 1224.395000 0.000000 1228.135000 0.630000 ;
      RECT 1219.715000 0.000000 1223.975000 0.630000 ;
      RECT 1215.140000 0.000000 1219.295000 0.630000 ;
      RECT 1210.560000 0.000000 1214.720000 0.630000 ;
      RECT 1205.985000 0.000000 1210.140000 0.630000 ;
      RECT 1201.410000 0.000000 1205.565000 0.630000 ;
      RECT 1196.730000 0.000000 1200.990000 0.630000 ;
      RECT 1192.155000 0.000000 1196.310000 0.630000 ;
      RECT 1187.995000 0.000000 1191.735000 0.630000 ;
      RECT 1183.420000 0.000000 1187.575000 0.630000 ;
      RECT 1178.840000 0.000000 1183.000000 0.630000 ;
      RECT 1174.160000 0.000000 1178.420000 0.630000 ;
      RECT 1169.585000 0.000000 1173.740000 0.630000 ;
      RECT 1165.115000 0.000000 1169.165000 0.630000 ;
      RECT 1160.540000 0.000000 1164.695000 0.630000 ;
      RECT 1155.960000 0.000000 1160.120000 0.630000 ;
      RECT 1151.800000 0.000000 1155.540000 0.630000 ;
      RECT 1147.225000 0.000000 1151.380000 0.630000 ;
      RECT 1142.650000 0.000000 1146.805000 0.630000 ;
      RECT 1138.075000 0.000000 1142.230000 0.630000 ;
      RECT 1133.500000 0.000000 1137.655000 0.630000 ;
      RECT 1128.820000 0.000000 1133.080000 0.630000 ;
      RECT 1124.240000 0.000000 1128.400000 0.630000 ;
      RECT 1119.770000 0.000000 1123.820000 0.630000 ;
      RECT 1115.610000 0.000000 1119.350000 0.630000 ;
      RECT 1110.825000 0.000000 1115.190000 0.630000 ;
      RECT 1106.355000 0.000000 1110.405000 0.630000 ;
      RECT 1101.780000 0.000000 1105.935000 0.630000 ;
      RECT 1097.200000 0.000000 1101.360000 0.630000 ;
      RECT 1092.625000 0.000000 1096.780000 0.630000 ;
      RECT 1087.945000 0.000000 1092.205000 0.630000 ;
      RECT 1083.370000 0.000000 1087.525000 0.630000 ;
      RECT 1079.210000 0.000000 1082.950000 0.630000 ;
      RECT 1074.635000 0.000000 1078.790000 0.630000 ;
      RECT 1070.060000 0.000000 1074.215000 0.630000 ;
      RECT 1065.380000 0.000000 1069.640000 0.630000 ;
      RECT 1060.800000 0.000000 1064.960000 0.630000 ;
      RECT 1056.225000 0.000000 1060.380000 0.630000 ;
      RECT 1051.755000 0.000000 1055.805000 0.630000 ;
      RECT 1047.180000 0.000000 1051.335000 0.630000 ;
      RECT 1042.810000 0.000000 1046.760000 0.630000 ;
      RECT 1038.340000 0.000000 1042.390000 0.630000 ;
      RECT 1033.760000 0.000000 1037.920000 0.630000 ;
      RECT 1029.185000 0.000000 1033.340000 0.630000 ;
      RECT 1024.505000 0.000000 1028.765000 0.630000 ;
      RECT 1019.930000 0.000000 1024.085000 0.630000 ;
      RECT 1015.355000 0.000000 1019.510000 0.630000 ;
      RECT 1010.780000 0.000000 1014.935000 0.630000 ;
      RECT 1006.200000 0.000000 1010.360000 0.630000 ;
      RECT 1002.040000 0.000000 1005.780000 0.630000 ;
      RECT 997.465000 0.000000 1001.620000 0.630000 ;
      RECT 992.995000 0.000000 997.045000 0.630000 ;
      RECT 988.420000 0.000000 992.575000 0.630000 ;
      RECT 983.840000 0.000000 988.000000 0.630000 ;
      RECT 979.160000 0.000000 983.420000 0.630000 ;
      RECT 974.585000 0.000000 978.740000 0.630000 ;
      RECT 970.010000 0.000000 974.165000 0.630000 ;
      RECT 965.850000 0.000000 969.590000 0.630000 ;
      RECT 961.275000 0.000000 965.430000 0.630000 ;
      RECT 956.700000 0.000000 960.855000 0.630000 ;
      RECT 952.020000 0.000000 956.280000 0.630000 ;
      RECT 947.440000 0.000000 951.600000 0.630000 ;
      RECT 942.865000 0.000000 947.020000 0.630000 ;
      RECT 938.290000 0.000000 942.445000 0.630000 ;
      RECT 933.610000 0.000000 937.870000 0.630000 ;
      RECT 929.450000 0.000000 933.190000 0.630000 ;
      RECT 924.875000 0.000000 929.030000 0.630000 ;
      RECT 920.400000 0.000000 924.455000 0.630000 ;
      RECT 915.620000 0.000000 919.980000 0.630000 ;
      RECT 911.145000 0.000000 915.200000 0.630000 ;
      RECT 906.570000 0.000000 910.725000 0.630000 ;
      RECT 901.995000 0.000000 906.150000 0.630000 ;
      RECT 897.420000 0.000000 901.575000 0.630000 ;
      RECT 893.260000 0.000000 897.000000 0.630000 ;
      RECT 888.680000 0.000000 892.840000 0.630000 ;
      RECT 884.105000 0.000000 888.260000 0.630000 ;
      RECT 879.530000 0.000000 883.685000 0.630000 ;
      RECT 875.060000 0.000000 879.110000 0.630000 ;
      RECT 870.275000 0.000000 874.640000 0.630000 ;
      RECT 865.800000 0.000000 869.855000 0.630000 ;
      RECT 861.225000 0.000000 865.380000 0.630000 ;
      RECT 857.065000 0.000000 860.805000 0.630000 ;
      RECT 852.385000 0.000000 856.645000 0.630000 ;
      RECT 847.810000 0.000000 851.965000 0.630000 ;
      RECT 843.235000 0.000000 847.390000 0.630000 ;
      RECT 838.660000 0.000000 842.815000 0.630000 ;
      RECT 834.080000 0.000000 838.240000 0.630000 ;
      RECT 829.400000 0.000000 833.660000 0.630000 ;
      RECT 824.825000 0.000000 828.980000 0.630000 ;
      RECT 820.665000 0.000000 824.405000 0.630000 ;
      RECT 816.090000 0.000000 820.245000 0.630000 ;
      RECT 811.515000 0.000000 815.670000 0.630000 ;
      RECT 807.040000 0.000000 811.095000 0.630000 ;
      RECT 802.260000 0.000000 806.620000 0.630000 ;
      RECT 797.785000 0.000000 801.840000 0.630000 ;
      RECT 793.210000 0.000000 797.365000 0.630000 ;
      RECT 788.635000 0.000000 792.790000 0.630000 ;
      RECT 784.475000 0.000000 788.215000 0.630000 ;
      RECT 779.900000 0.000000 784.055000 0.630000 ;
      RECT 775.320000 0.000000 779.480000 0.630000 ;
      RECT 770.745000 0.000000 774.900000 0.630000 ;
      RECT 766.170000 0.000000 770.325000 0.630000 ;
      RECT 761.490000 0.000000 765.750000 0.630000 ;
      RECT 756.915000 0.000000 761.070000 0.630000 ;
      RECT 752.440000 0.000000 756.495000 0.630000 ;
      RECT 748.280000 0.000000 752.020000 0.630000 ;
      RECT 743.500000 0.000000 747.860000 0.630000 ;
      RECT 739.025000 0.000000 743.080000 0.630000 ;
      RECT 734.450000 0.000000 738.605000 0.630000 ;
      RECT 729.875000 0.000000 734.030000 0.630000 ;
      RECT 725.300000 0.000000 729.455000 0.630000 ;
      RECT 720.620000 0.000000 724.880000 0.630000 ;
      RECT 716.040000 0.000000 720.200000 0.630000 ;
      RECT 711.880000 0.000000 715.620000 0.630000 ;
      RECT 707.305000 0.000000 711.460000 0.630000 ;
      RECT 702.730000 0.000000 706.885000 0.630000 ;
      RECT 698.155000 0.000000 702.310000 0.630000 ;
      RECT 693.475000 0.000000 697.735000 0.630000 ;
      RECT 688.900000 0.000000 693.055000 0.630000 ;
      RECT 684.425000 0.000000 688.480000 0.630000 ;
      RECT 679.850000 0.000000 684.005000 0.630000 ;
      RECT 675.690000 0.000000 679.430000 0.630000 ;
      RECT 671.010000 0.000000 675.270000 0.630000 ;
      RECT 666.435000 0.000000 670.590000 0.630000 ;
      RECT 661.860000 0.000000 666.015000 0.630000 ;
      RECT 657.280000 0.000000 661.440000 0.630000 ;
      RECT 652.600000 0.000000 656.860000 0.630000 ;
      RECT 648.025000 0.000000 652.180000 0.630000 ;
      RECT 643.450000 0.000000 647.605000 0.630000 ;
      RECT 639.395000 0.000000 643.030000 0.630000 ;
      RECT 634.715000 0.000000 638.975000 0.630000 ;
      RECT 630.140000 0.000000 634.295000 0.630000 ;
      RECT 625.665000 0.000000 629.720000 0.630000 ;
      RECT 621.090000 0.000000 625.245000 0.630000 ;
      RECT 616.515000 0.000000 620.670000 0.630000 ;
      RECT 611.835000 0.000000 616.095000 0.630000 ;
      RECT 607.260000 0.000000 611.415000 0.630000 ;
      RECT 603.200000 0.000000 606.840000 0.630000 ;
      RECT 598.520000 0.000000 602.780000 0.630000 ;
      RECT 593.945000 0.000000 598.100000 0.630000 ;
      RECT 589.370000 0.000000 593.525000 0.630000 ;
      RECT 584.795000 0.000000 588.950000 0.630000 ;
      RECT 580.115000 0.000000 584.375000 0.630000 ;
      RECT 575.540000 0.000000 579.695000 0.630000 ;
      RECT 570.960000 0.000000 575.120000 0.630000 ;
      RECT 566.800000 0.000000 570.540000 0.630000 ;
      RECT 562.120000 0.000000 566.380000 0.630000 ;
      RECT 557.545000 0.000000 561.700000 0.630000 ;
      RECT 553.075000 0.000000 557.125000 0.630000 ;
      RECT 548.500000 0.000000 552.655000 0.630000 ;
      RECT 543.820000 0.000000 548.080000 0.630000 ;
      RECT 539.240000 0.000000 543.400000 0.630000 ;
      RECT 534.665000 0.000000 538.820000 0.630000 ;
      RECT 530.610000 0.000000 534.245000 0.630000 ;
      RECT 525.930000 0.000000 530.190000 0.630000 ;
      RECT 521.355000 0.000000 525.510000 0.630000 ;
      RECT 516.780000 0.000000 520.935000 0.630000 ;
      RECT 512.200000 0.000000 516.360000 0.630000 ;
      RECT 507.730000 0.000000 511.780000 0.630000 ;
      RECT 502.945000 0.000000 507.310000 0.630000 ;
      RECT 498.475000 0.000000 502.525000 0.630000 ;
      RECT 493.900000 0.000000 498.055000 0.630000 ;
      RECT 489.740000 0.000000 493.480000 0.630000 ;
      RECT 485.060000 0.000000 489.320000 0.630000 ;
      RECT 480.480000 0.000000 484.640000 0.630000 ;
      RECT 475.905000 0.000000 480.060000 0.630000 ;
      RECT 471.330000 0.000000 475.485000 0.630000 ;
      RECT 466.755000 0.000000 470.910000 0.630000 ;
      RECT 462.075000 0.000000 466.335000 0.630000 ;
      RECT 457.500000 0.000000 461.655000 0.630000 ;
      RECT 453.440000 0.000000 457.080000 0.630000 ;
      RECT 448.760000 0.000000 453.020000 0.630000 ;
      RECT 444.185000 0.000000 448.340000 0.630000 ;
      RECT 439.715000 0.000000 443.765000 0.630000 ;
      RECT 435.140000 0.000000 439.295000 0.630000 ;
      RECT 430.460000 0.000000 434.720000 0.630000 ;
      RECT 425.880000 0.000000 430.040000 0.630000 ;
      RECT 421.305000 0.000000 425.460000 0.630000 ;
      RECT 417.145000 0.000000 420.885000 0.630000 ;
      RECT 412.570000 0.000000 416.725000 0.630000 ;
      RECT 407.995000 0.000000 412.150000 0.630000 ;
      RECT 403.420000 0.000000 407.575000 0.630000 ;
      RECT 398.840000 0.000000 403.000000 0.630000 ;
      RECT 394.160000 0.000000 398.420000 0.630000 ;
      RECT 389.585000 0.000000 393.740000 0.630000 ;
      RECT 385.115000 0.000000 389.165000 0.630000 ;
      RECT 380.955000 0.000000 384.695000 0.630000 ;
      RECT 376.170000 0.000000 380.535000 0.630000 ;
      RECT 371.700000 0.000000 375.750000 0.630000 ;
      RECT 367.120000 0.000000 371.280000 0.630000 ;
      RECT 362.545000 0.000000 366.700000 0.630000 ;
      RECT 357.970000 0.000000 362.125000 0.630000 ;
      RECT 353.290000 0.000000 357.550000 0.630000 ;
      RECT 348.715000 0.000000 352.870000 0.630000 ;
      RECT 344.660000 0.000000 348.295000 0.630000 ;
      RECT 339.980000 0.000000 344.240000 0.630000 ;
      RECT 335.400000 0.000000 339.560000 0.630000 ;
      RECT 330.825000 0.000000 334.980000 0.630000 ;
      RECT 326.355000 0.000000 330.405000 0.630000 ;
      RECT 321.570000 0.000000 325.935000 0.630000 ;
      RECT 317.100000 0.000000 321.150000 0.630000 ;
      RECT 312.520000 0.000000 316.680000 0.630000 ;
      RECT 308.360000 0.000000 312.100000 0.630000 ;
      RECT 303.785000 0.000000 307.940000 0.630000 ;
      RECT 299.105000 0.000000 303.365000 0.630000 ;
      RECT 294.530000 0.000000 298.685000 0.630000 ;
      RECT 289.955000 0.000000 294.110000 0.630000 ;
      RECT 285.380000 0.000000 289.535000 0.630000 ;
      RECT 280.700000 0.000000 284.960000 0.630000 ;
      RECT 276.120000 0.000000 280.280000 0.630000 ;
      RECT 272.065000 0.000000 275.700000 0.630000 ;
      RECT 267.385000 0.000000 271.645000 0.630000 ;
      RECT 262.810000 0.000000 266.965000 0.630000 ;
      RECT 258.235000 0.000000 262.390000 0.630000 ;
      RECT 253.760000 0.000000 257.815000 0.630000 ;
      RECT 249.185000 0.000000 253.340000 0.630000 ;
      RECT 244.505000 0.000000 248.765000 0.630000 ;
      RECT 239.930000 0.000000 244.085000 0.630000 ;
      RECT 235.875000 0.000000 239.510000 0.630000 ;
      RECT 231.300000 0.000000 235.455000 0.630000 ;
      RECT 226.620000 0.000000 230.880000 0.630000 ;
      RECT 222.040000 0.000000 226.200000 0.630000 ;
      RECT 217.465000 0.000000 221.620000 0.630000 ;
      RECT 212.785000 0.000000 217.045000 0.630000 ;
      RECT 208.210000 0.000000 212.365000 0.630000 ;
      RECT 203.635000 0.000000 207.790000 0.630000 ;
      RECT 199.475000 0.000000 203.215000 0.630000 ;
      RECT 195.000000 0.000000 199.055000 0.630000 ;
      RECT 190.220000 0.000000 194.580000 0.630000 ;
      RECT 185.745000 0.000000 189.800000 0.630000 ;
      RECT 181.170000 0.000000 185.325000 0.630000 ;
      RECT 176.595000 0.000000 180.750000 0.630000 ;
      RECT 171.915000 0.000000 176.175000 0.630000 ;
      RECT 167.340000 0.000000 171.495000 0.630000 ;
      RECT 163.280000 0.000000 166.920000 0.630000 ;
      RECT 158.600000 0.000000 162.860000 0.630000 ;
      RECT 154.025000 0.000000 158.180000 0.630000 ;
      RECT 149.450000 0.000000 153.605000 0.630000 ;
      RECT 144.875000 0.000000 149.030000 0.630000 ;
      RECT 140.400000 0.000000 144.455000 0.630000 ;
      RECT 135.620000 0.000000 139.980000 0.630000 ;
      RECT 131.145000 0.000000 135.200000 0.630000 ;
      RECT 126.985000 0.000000 130.725000 0.630000 ;
      RECT 122.410000 0.000000 126.565000 0.630000 ;
      RECT 117.730000 0.000000 121.990000 0.630000 ;
      RECT 113.155000 0.000000 117.310000 0.630000 ;
      RECT 108.580000 0.000000 112.735000 0.630000 ;
      RECT 104.000000 0.000000 108.160000 0.630000 ;
      RECT 99.425000 0.000000 103.580000 0.630000 ;
      RECT 94.745000 0.000000 99.005000 0.630000 ;
      RECT 90.690000 0.000000 94.325000 0.630000 ;
      RECT 86.115000 0.000000 90.270000 0.630000 ;
      RECT 81.640000 0.000000 85.695000 0.630000 ;
      RECT 76.860000 0.000000 81.220000 0.630000 ;
      RECT 72.385000 0.000000 76.440000 0.630000 ;
      RECT 67.810000 0.000000 71.965000 0.630000 ;
      RECT 63.130000 0.000000 67.390000 0.630000 ;
      RECT 58.555000 0.000000 62.710000 0.630000 ;
      RECT 54.500000 0.000000 58.135000 0.630000 ;
      RECT 49.820000 0.000000 54.080000 0.630000 ;
      RECT 45.240000 0.000000 49.400000 0.630000 ;
      RECT 40.665000 0.000000 44.820000 0.630000 ;
      RECT 36.090000 0.000000 40.245000 0.630000 ;
      RECT 31.515000 0.000000 35.670000 0.630000 ;
      RECT 26.835000 0.000000 31.095000 0.630000 ;
      RECT 22.260000 0.000000 26.415000 0.630000 ;
      RECT 18.100000 0.000000 21.840000 0.630000 ;
      RECT 13.625000 0.000000 17.680000 0.630000 ;
      RECT 8.840000 0.000000 13.205000 0.630000 ;
      RECT 6.660000 0.000000 8.420000 0.625000 ;
      RECT 4.370000 0.000000 6.240000 0.625000 ;
      RECT 0.000000 0.000000 3.950000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 2056.950000 2299.540000 2118.880000 ;
      RECT 1.100000 2056.250000 2299.540000 2056.950000 ;
      RECT 1.100000 2056.050000 2298.440000 2056.250000 ;
      RECT 0.000000 2055.350000 2298.440000 2056.050000 ;
      RECT 0.000000 2021.550000 2299.540000 2055.350000 ;
      RECT 1.100000 2020.650000 2299.540000 2021.550000 ;
      RECT 0.000000 2020.150000 2299.540000 2020.650000 ;
      RECT 0.000000 2019.250000 2298.440000 2020.150000 ;
      RECT 0.000000 1982.750000 2299.540000 2019.250000 ;
      RECT 1.100000 1981.850000 2299.540000 1982.750000 ;
      RECT 0.000000 1980.550000 2299.540000 1981.850000 ;
      RECT 0.000000 1979.650000 2298.440000 1980.550000 ;
      RECT 0.000000 1943.750000 2299.540000 1979.650000 ;
      RECT 1.100000 1942.850000 2299.540000 1943.750000 ;
      RECT 0.000000 1941.150000 2299.540000 1942.850000 ;
      RECT 0.000000 1940.250000 2298.440000 1941.150000 ;
      RECT 0.000000 1905.050000 2299.540000 1940.250000 ;
      RECT 1.100000 1904.150000 2299.540000 1905.050000 ;
      RECT 0.000000 1901.650000 2299.540000 1904.150000 ;
      RECT 0.000000 1900.750000 2298.440000 1901.650000 ;
      RECT 0.000000 1866.050000 2299.540000 1900.750000 ;
      RECT 1.100000 1865.150000 2299.540000 1866.050000 ;
      RECT 0.000000 1861.850000 2299.540000 1865.150000 ;
      RECT 0.000000 1860.950000 2298.440000 1861.850000 ;
      RECT 0.000000 1827.050000 2299.540000 1860.950000 ;
      RECT 1.100000 1826.150000 2299.540000 1827.050000 ;
      RECT 0.000000 1822.350000 2299.540000 1826.150000 ;
      RECT 0.000000 1821.450000 2298.440000 1822.350000 ;
      RECT 0.000000 1788.450000 2299.540000 1821.450000 ;
      RECT 1.100000 1787.550000 2299.540000 1788.450000 ;
      RECT 0.000000 1782.750000 2299.540000 1787.550000 ;
      RECT 0.000000 1781.850000 2298.440000 1782.750000 ;
      RECT 0.000000 1749.350000 2299.540000 1781.850000 ;
      RECT 1.100000 1748.450000 2299.540000 1749.350000 ;
      RECT 0.000000 1742.950000 2299.540000 1748.450000 ;
      RECT 0.000000 1742.050000 2298.440000 1742.950000 ;
      RECT 0.000000 1710.650000 2299.540000 1742.050000 ;
      RECT 1.100000 1709.750000 2299.540000 1710.650000 ;
      RECT 0.000000 1703.450000 2299.540000 1709.750000 ;
      RECT 0.000000 1702.550000 2298.440000 1703.450000 ;
      RECT 0.000000 1671.550000 2299.540000 1702.550000 ;
      RECT 1.100000 1670.650000 2299.540000 1671.550000 ;
      RECT 0.000000 1663.950000 2299.540000 1670.650000 ;
      RECT 0.000000 1663.050000 2298.440000 1663.950000 ;
      RECT 0.000000 1632.950000 2299.540000 1663.050000 ;
      RECT 1.100000 1632.050000 2299.540000 1632.950000 ;
      RECT 0.000000 1624.050000 2299.540000 1632.050000 ;
      RECT 0.000000 1623.150000 2298.440000 1624.050000 ;
      RECT 0.000000 1594.050000 2299.540000 1623.150000 ;
      RECT 1.100000 1593.150000 2299.540000 1594.050000 ;
      RECT 0.000000 1584.650000 2299.540000 1593.150000 ;
      RECT 0.000000 1583.750000 2298.440000 1584.650000 ;
      RECT 0.000000 1555.250000 2299.540000 1583.750000 ;
      RECT 1.100000 1554.350000 2299.540000 1555.250000 ;
      RECT 0.000000 1545.150000 2299.540000 1554.350000 ;
      RECT 0.000000 1544.250000 2298.440000 1545.150000 ;
      RECT 0.000000 1516.350000 2299.540000 1544.250000 ;
      RECT 1.100000 1515.450000 2299.540000 1516.350000 ;
      RECT 0.000000 1505.250000 2299.540000 1515.450000 ;
      RECT 0.000000 1504.350000 2298.440000 1505.250000 ;
      RECT 0.000000 1477.150000 2299.540000 1504.350000 ;
      RECT 1.100000 1476.250000 2299.540000 1477.150000 ;
      RECT 0.000000 1465.650000 2299.540000 1476.250000 ;
      RECT 0.000000 1464.750000 2298.440000 1465.650000 ;
      RECT 0.000000 1438.550000 2299.540000 1464.750000 ;
      RECT 1.100000 1437.650000 2299.540000 1438.550000 ;
      RECT 0.000000 1426.250000 2299.540000 1437.650000 ;
      RECT 0.000000 1425.350000 2298.440000 1426.250000 ;
      RECT 0.000000 1399.350000 2299.540000 1425.350000 ;
      RECT 1.100000 1398.450000 2299.540000 1399.350000 ;
      RECT 0.000000 1386.250000 2299.540000 1398.450000 ;
      RECT 0.000000 1385.350000 2298.440000 1386.250000 ;
      RECT 0.000000 1360.950000 2299.540000 1385.350000 ;
      RECT 1.100000 1360.050000 2299.540000 1360.950000 ;
      RECT 0.000000 1346.850000 2299.540000 1360.050000 ;
      RECT 0.000000 1345.950000 2298.440000 1346.850000 ;
      RECT 0.000000 1321.850000 2299.540000 1345.950000 ;
      RECT 1.100000 1320.950000 2299.540000 1321.850000 ;
      RECT 0.000000 1307.350000 2299.540000 1320.950000 ;
      RECT 0.000000 1306.450000 2298.440000 1307.350000 ;
      RECT 0.000000 1283.150000 2299.540000 1306.450000 ;
      RECT 1.100000 1282.250000 2299.540000 1283.150000 ;
      RECT 0.000000 1267.450000 2299.540000 1282.250000 ;
      RECT 0.000000 1266.550000 2298.440000 1267.450000 ;
      RECT 0.000000 1244.150000 2299.540000 1266.550000 ;
      RECT 1.100000 1243.250000 2299.540000 1244.150000 ;
      RECT 0.000000 1227.950000 2299.540000 1243.250000 ;
      RECT 0.000000 1227.050000 2298.440000 1227.950000 ;
      RECT 0.000000 1205.450000 2299.540000 1227.050000 ;
      RECT 1.100000 1204.550000 2299.540000 1205.450000 ;
      RECT 0.000000 1188.450000 2299.540000 1204.550000 ;
      RECT 0.000000 1187.550000 2298.440000 1188.450000 ;
      RECT 0.000000 1166.350000 2299.540000 1187.550000 ;
      RECT 1.100000 1165.450000 2299.540000 1166.350000 ;
      RECT 0.000000 1149.050000 2299.540000 1165.450000 ;
      RECT 0.000000 1148.150000 2298.440000 1149.050000 ;
      RECT 0.000000 1127.350000 2299.540000 1148.150000 ;
      RECT 1.100000 1126.450000 2299.540000 1127.350000 ;
      RECT 0.000000 1109.150000 2299.540000 1126.450000 ;
      RECT 0.000000 1108.250000 2298.440000 1109.150000 ;
      RECT 0.000000 1088.850000 2299.540000 1108.250000 ;
      RECT 1.100000 1087.950000 2299.540000 1088.850000 ;
      RECT 0.000000 1069.650000 2299.540000 1087.950000 ;
      RECT 0.000000 1068.750000 2298.440000 1069.650000 ;
      RECT 0.000000 1049.650000 2299.540000 1068.750000 ;
      RECT 1.100000 1048.750000 2299.540000 1049.650000 ;
      RECT 0.000000 1030.150000 2299.540000 1048.750000 ;
      RECT 0.000000 1029.250000 2298.440000 1030.150000 ;
      RECT 0.000000 1011.150000 2299.540000 1029.250000 ;
      RECT 1.100000 1010.250000 2299.540000 1011.150000 ;
      RECT 0.000000 990.350000 2299.540000 1010.250000 ;
      RECT 0.000000 989.450000 2298.440000 990.350000 ;
      RECT 0.000000 971.850000 2299.540000 989.450000 ;
      RECT 1.100000 970.950000 2299.540000 971.850000 ;
      RECT 0.000000 950.650000 2299.540000 970.950000 ;
      RECT 0.000000 949.750000 2298.440000 950.650000 ;
      RECT 0.000000 933.350000 2299.540000 949.750000 ;
      RECT 1.100000 932.450000 2299.540000 933.350000 ;
      RECT 0.000000 911.250000 2299.540000 932.450000 ;
      RECT 0.000000 910.350000 2298.440000 911.250000 ;
      RECT 0.000000 894.350000 2299.540000 910.350000 ;
      RECT 1.100000 893.450000 2299.540000 894.350000 ;
      RECT 0.000000 871.350000 2299.540000 893.450000 ;
      RECT 0.000000 870.450000 2298.440000 871.350000 ;
      RECT 0.000000 855.650000 2299.540000 870.450000 ;
      RECT 1.100000 854.750000 2299.540000 855.650000 ;
      RECT 0.000000 831.950000 2299.540000 854.750000 ;
      RECT 0.000000 831.050000 2298.440000 831.950000 ;
      RECT 0.000000 816.650000 2299.540000 831.050000 ;
      RECT 1.100000 815.750000 2299.540000 816.650000 ;
      RECT 0.000000 792.450000 2299.540000 815.750000 ;
      RECT 0.000000 791.550000 2298.440000 792.450000 ;
      RECT 0.000000 777.550000 2299.540000 791.550000 ;
      RECT 1.100000 776.650000 2299.540000 777.550000 ;
      RECT 0.000000 752.550000 2299.540000 776.650000 ;
      RECT 0.000000 751.650000 2298.440000 752.550000 ;
      RECT 0.000000 739.050000 2299.540000 751.650000 ;
      RECT 1.100000 738.150000 2299.540000 739.050000 ;
      RECT 0.000000 713.050000 2299.540000 738.150000 ;
      RECT 0.000000 712.150000 2298.440000 713.050000 ;
      RECT 0.000000 699.850000 2299.540000 712.150000 ;
      RECT 1.100000 698.950000 2299.540000 699.850000 ;
      RECT 0.000000 673.550000 2299.540000 698.950000 ;
      RECT 0.000000 672.650000 2298.440000 673.550000 ;
      RECT 0.000000 661.350000 2299.540000 672.650000 ;
      RECT 1.100000 660.450000 2299.540000 661.350000 ;
      RECT 0.000000 633.650000 2299.540000 660.450000 ;
      RECT 0.000000 632.750000 2298.440000 633.650000 ;
      RECT 0.000000 622.150000 2299.540000 632.750000 ;
      RECT 1.100000 621.250000 2299.540000 622.150000 ;
      RECT 0.000000 594.150000 2299.540000 621.250000 ;
      RECT 0.000000 593.250000 2298.440000 594.150000 ;
      RECT 0.000000 583.650000 2299.540000 593.250000 ;
      RECT 1.100000 582.750000 2299.540000 583.650000 ;
      RECT 0.000000 554.750000 2299.540000 582.750000 ;
      RECT 0.000000 553.850000 2298.440000 554.750000 ;
      RECT 0.000000 544.550000 2299.540000 553.850000 ;
      RECT 1.100000 543.650000 2299.540000 544.550000 ;
      RECT 0.000000 514.850000 2299.540000 543.650000 ;
      RECT 0.000000 513.950000 2298.440000 514.850000 ;
      RECT 0.000000 505.950000 2299.540000 513.950000 ;
      RECT 1.100000 505.050000 2299.540000 505.950000 ;
      RECT 0.000000 475.350000 2299.540000 505.050000 ;
      RECT 0.000000 474.450000 2298.440000 475.350000 ;
      RECT 0.000000 466.750000 2299.540000 474.450000 ;
      RECT 1.100000 465.850000 2299.540000 466.750000 ;
      RECT 0.000000 435.750000 2299.540000 465.850000 ;
      RECT 0.000000 434.850000 2298.440000 435.750000 ;
      RECT 0.000000 427.850000 2299.540000 434.850000 ;
      RECT 1.100000 426.950000 2299.540000 427.850000 ;
      RECT 0.000000 396.350000 2299.540000 426.950000 ;
      RECT 0.000000 395.450000 2298.440000 396.350000 ;
      RECT 0.000000 389.150000 2299.540000 395.450000 ;
      RECT 1.100000 388.250000 2299.540000 389.150000 ;
      RECT 0.000000 356.350000 2299.540000 388.250000 ;
      RECT 0.000000 355.450000 2298.440000 356.350000 ;
      RECT 0.000000 350.050000 2299.540000 355.450000 ;
      RECT 1.100000 349.150000 2299.540000 350.050000 ;
      RECT 0.000000 317.050000 2299.540000 349.150000 ;
      RECT 0.000000 316.150000 2298.440000 317.050000 ;
      RECT 0.000000 311.550000 2299.540000 316.150000 ;
      RECT 1.100000 310.650000 2299.540000 311.550000 ;
      RECT 0.000000 277.550000 2299.540000 310.650000 ;
      RECT 0.000000 276.650000 2298.440000 277.550000 ;
      RECT 0.000000 272.350000 2299.540000 276.650000 ;
      RECT 1.100000 271.450000 2299.540000 272.350000 ;
      RECT 0.000000 237.550000 2299.540000 271.450000 ;
      RECT 0.000000 236.650000 2298.440000 237.550000 ;
      RECT 0.000000 233.850000 2299.540000 236.650000 ;
      RECT 1.100000 232.950000 2299.540000 233.850000 ;
      RECT 0.000000 198.050000 2299.540000 232.950000 ;
      RECT 0.000000 197.150000 2298.440000 198.050000 ;
      RECT 0.000000 194.650000 2299.540000 197.150000 ;
      RECT 1.100000 193.750000 2299.540000 194.650000 ;
      RECT 0.000000 158.650000 2299.540000 193.750000 ;
      RECT 0.000000 157.750000 2298.440000 158.650000 ;
      RECT 0.000000 156.150000 2299.540000 157.750000 ;
      RECT 1.100000 155.250000 2299.540000 156.150000 ;
      RECT 0.000000 118.650000 2299.540000 155.250000 ;
      RECT 0.000000 117.750000 2298.440000 118.650000 ;
      RECT 0.000000 117.050000 2299.540000 117.750000 ;
      RECT 1.100000 116.150000 2299.540000 117.050000 ;
      RECT 0.000000 79.250000 2299.540000 116.150000 ;
      RECT 0.000000 78.350000 2298.440000 79.250000 ;
      RECT 0.000000 78.050000 2299.540000 78.350000 ;
      RECT 1.100000 77.150000 2299.540000 78.050000 ;
      RECT 0.000000 39.850000 2299.540000 77.150000 ;
      RECT 0.000000 39.350000 2298.440000 39.850000 ;
      RECT 1.100000 38.950000 2298.440000 39.350000 ;
      RECT 1.100000 38.450000 2299.540000 38.950000 ;
      RECT 0.000000 4.150000 2299.540000 38.450000 ;
      RECT 1.100000 3.350000 2299.540000 4.150000 ;
      RECT 1.100000 3.250000 2298.440000 3.350000 ;
      RECT 0.000000 2.450000 2298.440000 3.250000 ;
      RECT 0.000000 0.000000 2299.540000 2.450000 ;
    LAYER met4 ;
      RECT 0.000000 2104.800000 2299.540000 2118.880000 ;
      RECT 23.420000 2092.800000 2276.120000 2104.800000 ;
      RECT 2274.920000 24.720000 2276.120000 2092.800000 ;
      RECT 35.420000 24.720000 2264.120000 2092.800000 ;
      RECT 23.420000 24.720000 24.620000 2092.800000 ;
      RECT 2286.920000 12.720000 2299.540000 2104.800000 ;
      RECT 23.420000 12.720000 2276.120000 24.720000 ;
      RECT 0.000000 12.720000 12.620000 2104.800000 ;
      RECT 0.000000 0.000000 2299.540000 12.720000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
