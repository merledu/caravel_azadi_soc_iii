##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Thu Mar 17 14:21:38 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2369.460000 BY 2290.240000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.430000 0.000000 4.570000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.530000 0.000000 1.670000 0.490000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.230000 0.000000 468.370000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.530000 0.000000 157.670000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.730000 0.000000 472.870000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.730000 0.000000 463.870000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.230000 0.000000 459.370000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.730000 0.000000 454.870000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.230000 0.000000 450.370000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.630000 0.000000 301.770000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.130000 0.000000 297.270000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.530000 0.000000 292.670000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.030000 0.000000 288.170000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.530000 0.000000 283.670000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.030000 0.000000 279.170000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.530000 0.000000 274.670000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.030000 0.000000 270.170000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.530000 0.000000 265.670000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.030000 0.000000 261.170000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.530000 0.000000 256.670000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.030000 0.000000 252.170000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.530000 0.000000 247.670000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.030000 0.000000 243.170000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.530000 0.000000 238.670000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.030000 0.000000 234.170000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.530000 0.000000 229.670000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030000 0.000000 225.170000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.530000 0.000000 220.670000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.030000 0.000000 216.170000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.530000 0.000000 211.670000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.030000 0.000000 207.170000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.530000 0.000000 202.670000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.030000 0.000000 198.170000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.530000 0.000000 193.670000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.030000 0.000000 189.170000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.530000 0.000000 184.670000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.030000 0.000000 180.170000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.530000 0.000000 175.670000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.030000 0.000000 171.170000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.530000 0.000000 166.670000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.030000 0.000000 162.170000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.030000 0.000000 153.170000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.530000 0.000000 148.670000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.930000 0.000000 144.070000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.430000 0.000000 139.570000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.930000 0.000000 135.070000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.430000 0.000000 130.570000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.930000 0.000000 126.070000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.430000 0.000000 121.570000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930000 0.000000 117.070000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.430000 0.000000 112.570000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.930000 0.000000 108.070000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.430000 0.000000 103.570000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.930000 0.000000 99.070000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.430000 0.000000 94.570000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.930000 0.000000 90.070000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.430000 0.000000 85.570000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.930000 0.000000 81.070000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.430000 0.000000 76.570000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.930000 0.000000 72.070000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.430000 0.000000 67.570000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.930000 0.000000 63.070000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.430000 0.000000 58.570000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.930000 0.000000 54.070000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.430000 0.000000 49.570000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.930000 0.000000 45.070000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430000 0.000000 40.570000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.930000 0.000000 36.070000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.430000 0.000000 31.570000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.930000 0.000000 27.070000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.430000 0.000000 22.570000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.930000 0.000000 18.070000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430000 0.000000 13.570000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.930000 0.000000 9.070000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.630000 0.000000 445.770000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.130000 0.000000 441.270000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630000 0.000000 436.770000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.130000 0.000000 432.270000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.630000 0.000000 427.770000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.130000 0.000000 423.270000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.630000 0.000000 418.770000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.130000 0.000000 414.270000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.630000 0.000000 409.770000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.130000 0.000000 405.270000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.630000 0.000000 400.770000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.130000 0.000000 396.270000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.630000 0.000000 391.770000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.130000 0.000000 387.270000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.630000 0.000000 382.770000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.130000 0.000000 378.270000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.630000 0.000000 373.770000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.130000 0.000000 369.270000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.630000 0.000000 364.770000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.130000 0.000000 360.270000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.630000 0.000000 355.770000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.130000 0.000000 351.270000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.630000 0.000000 346.770000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.130000 0.000000 342.270000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.630000 0.000000 337.770000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130000 0.000000 333.270000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.630000 0.000000 328.770000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.130000 0.000000 324.270000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.630000 0.000000 319.770000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.130000 0.000000 315.270000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.630000 0.000000 310.770000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.130000 0.000000 306.270000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.130000 0.000000 1049.270000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.530000 0.000000 1044.670000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.030000 0.000000 1040.170000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.530000 0.000000 1035.670000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.030000 0.000000 1031.170000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.530000 0.000000 1026.670000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.030000 0.000000 1022.170000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.530000 0.000000 1017.670000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.030000 0.000000 1013.170000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.530000 0.000000 1008.670000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.030000 0.000000 1004.170000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.530000 0.000000 999.670000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.030000 0.000000 995.170000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.530000 0.000000 990.670000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.030000 0.000000 986.170000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.530000 0.000000 981.670000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.030000 0.000000 977.170000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530000 0.000000 972.670000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.030000 0.000000 968.170000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.530000 0.000000 963.670000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.030000 0.000000 959.170000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.530000 0.000000 954.670000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.030000 0.000000 950.170000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.530000 0.000000 945.670000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.030000 0.000000 941.170000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.530000 0.000000 936.670000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.030000 0.000000 932.170000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.530000 0.000000 927.670000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.030000 0.000000 923.170000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.530000 0.000000 918.670000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.030000 0.000000 914.170000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.530000 0.000000 909.670000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.030000 0.000000 905.170000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.530000 0.000000 900.670000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.930000 0.000000 896.070000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.430000 0.000000 891.570000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.930000 0.000000 887.070000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.430000 0.000000 882.570000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.930000 0.000000 878.070000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.430000 0.000000 873.570000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.930000 0.000000 869.070000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430000 0.000000 864.570000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.930000 0.000000 860.070000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.430000 0.000000 855.570000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.930000 0.000000 851.070000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.430000 0.000000 846.570000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.930000 0.000000 842.070000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.430000 0.000000 837.570000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.930000 0.000000 833.070000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.430000 0.000000 828.570000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.930000 0.000000 824.070000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.430000 0.000000 819.570000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.930000 0.000000 815.070000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.430000 0.000000 810.570000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.930000 0.000000 806.070000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.430000 0.000000 801.570000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.930000 0.000000 797.070000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.430000 0.000000 792.570000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.930000 0.000000 788.070000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.430000 0.000000 783.570000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.930000 0.000000 779.070000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.430000 0.000000 774.570000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.930000 0.000000 770.070000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.430000 0.000000 765.570000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930000 0.000000 761.070000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.430000 0.000000 756.570000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.930000 0.000000 752.070000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.430000 0.000000 747.570000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.830000 0.000000 742.970000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.330000 0.000000 738.470000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.830000 0.000000 733.970000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.330000 0.000000 729.470000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.830000 0.000000 724.970000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.330000 0.000000 720.470000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.830000 0.000000 715.970000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.330000 0.000000 711.470000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.830000 0.000000 706.970000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.330000 0.000000 702.470000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.830000 0.000000 697.970000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.330000 0.000000 693.470000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.830000 0.000000 688.970000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.330000 0.000000 684.470000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.830000 0.000000 679.970000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.330000 0.000000 675.470000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.830000 0.000000 670.970000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.330000 0.000000 666.470000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.830000 0.000000 661.970000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.330000 0.000000 657.470000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830000 0.000000 652.970000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.330000 0.000000 648.470000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.830000 0.000000 643.970000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.330000 0.000000 639.470000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.830000 0.000000 634.970000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.330000 0.000000 630.470000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.830000 0.000000 625.970000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.330000 0.000000 621.470000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.830000 0.000000 616.970000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.330000 0.000000 612.470000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.830000 0.000000 607.970000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.330000 0.000000 603.470000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.830000 0.000000 598.970000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.230000 0.000000 594.370000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.730000 0.000000 589.870000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.230000 0.000000 585.370000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.730000 0.000000 580.870000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.230000 0.000000 576.370000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.730000 0.000000 571.870000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.230000 0.000000 567.370000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.730000 0.000000 562.870000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.230000 0.000000 558.370000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.730000 0.000000 553.870000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.230000 0.000000 549.370000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730000 0.000000 544.870000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.230000 0.000000 540.370000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.730000 0.000000 535.870000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.230000 0.000000 531.370000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.730000 0.000000 526.870000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.230000 0.000000 522.370000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.730000 0.000000 517.870000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.230000 0.000000 513.370000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.730000 0.000000 508.870000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.230000 0.000000 504.370000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.730000 0.000000 499.870000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.230000 0.000000 495.370000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.730000 0.000000 490.870000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.230000 0.000000 486.370000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.730000 0.000000 481.870000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.230000 0.000000 477.370000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.430000 0.000000 1625.570000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.930000 0.000000 1621.070000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.430000 0.000000 1616.570000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.930000 0.000000 1612.070000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.430000 0.000000 1607.570000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.930000 0.000000 1603.070000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.430000 0.000000 1598.570000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.930000 0.000000 1594.070000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.430000 0.000000 1589.570000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.930000 0.000000 1585.070000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.430000 0.000000 1580.570000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.930000 0.000000 1576.070000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.430000 0.000000 1571.570000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.930000 0.000000 1567.070000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.430000 0.000000 1562.570000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.930000 0.000000 1558.070000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.430000 0.000000 1553.570000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.930000 0.000000 1549.070000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.430000 0.000000 1544.570000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.930000 0.000000 1540.070000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.430000 0.000000 1535.570000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.930000 0.000000 1531.070000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.430000 0.000000 1526.570000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.930000 0.000000 1522.070000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.430000 0.000000 1517.570000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.930000 0.000000 1513.070000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430000 0.000000 1508.570000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.930000 0.000000 1504.070000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.430000 0.000000 1499.570000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.830000 0.000000 1494.970000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.330000 0.000000 1490.470000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.830000 0.000000 1485.970000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.330000 0.000000 1481.470000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.830000 0.000000 1476.970000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.330000 0.000000 1472.470000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.830000 0.000000 1467.970000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.330000 0.000000 1463.470000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.830000 0.000000 1458.970000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.330000 0.000000 1454.470000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.830000 0.000000 1449.970000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.330000 0.000000 1445.470000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.830000 0.000000 1440.970000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.330000 0.000000 1436.470000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.830000 0.000000 1431.970000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.330000 0.000000 1427.470000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.830000 0.000000 1422.970000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.330000 0.000000 1418.470000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.830000 0.000000 1413.970000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.330000 0.000000 1409.470000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.830000 0.000000 1404.970000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.330000 0.000000 1400.470000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.830000 0.000000 1395.970000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.330000 0.000000 1391.470000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.830000 0.000000 1386.970000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.330000 0.000000 1382.470000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.830000 0.000000 1377.970000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.330000 0.000000 1373.470000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.830000 0.000000 1368.970000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.330000 0.000000 1364.470000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.830000 0.000000 1359.970000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.330000 0.000000 1355.470000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.830000 0.000000 1350.970000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.230000 0.000000 1346.370000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.730000 0.000000 1341.870000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.230000 0.000000 1337.370000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.730000 0.000000 1332.870000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.230000 0.000000 1328.370000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.730000 0.000000 1323.870000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.230000 0.000000 1319.370000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.730000 0.000000 1314.870000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.230000 0.000000 1310.370000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.730000 0.000000 1305.870000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.230000 0.000000 1301.370000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.730000 0.000000 1296.870000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.230000 0.000000 1292.370000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.730000 0.000000 1287.870000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.230000 0.000000 1283.370000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.730000 0.000000 1278.870000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.230000 0.000000 1274.370000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.730000 0.000000 1269.870000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.230000 0.000000 1265.370000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.730000 0.000000 1260.870000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.230000 0.000000 1256.370000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.730000 0.000000 1251.870000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.230000 0.000000 1247.370000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.730000 0.000000 1242.870000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.230000 0.000000 1238.370000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.730000 0.000000 1233.870000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.230000 0.000000 1229.370000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.730000 0.000000 1224.870000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.230000 0.000000 1220.370000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.730000 0.000000 1215.870000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.230000 0.000000 1211.370000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.730000 0.000000 1206.870000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.230000 0.000000 1202.370000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.730000 0.000000 1197.870000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.130000 0.000000 1193.270000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.630000 0.000000 1188.770000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130000 0.000000 1184.270000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.630000 0.000000 1179.770000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.130000 0.000000 1175.270000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.630000 0.000000 1170.770000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.130000 0.000000 1166.270000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.630000 0.000000 1161.770000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.130000 0.000000 1157.270000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.630000 0.000000 1152.770000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.130000 0.000000 1148.270000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.630000 0.000000 1143.770000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.130000 0.000000 1139.270000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.630000 0.000000 1134.770000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.130000 0.000000 1130.270000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.630000 0.000000 1125.770000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.130000 0.000000 1121.270000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.630000 0.000000 1116.770000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.130000 0.000000 1112.270000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630000 0.000000 1107.770000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.130000 0.000000 1103.270000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.630000 0.000000 1098.770000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.130000 0.000000 1094.270000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.630000 0.000000 1089.770000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.130000 0.000000 1085.270000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630000 0.000000 1080.770000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.130000 0.000000 1076.270000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.630000 0.000000 1071.770000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.130000 0.000000 1067.270000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.630000 0.000000 1062.770000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.130000 0.000000 1058.270000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.630000 0.000000 1053.770000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.830000 0.000000 2201.970000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.330000 0.000000 2197.470000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.830000 0.000000 2192.970000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.330000 0.000000 2188.470000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.830000 0.000000 2183.970000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.330000 0.000000 2179.470000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.830000 0.000000 2174.970000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.330000 0.000000 2170.470000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.830000 0.000000 2165.970000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.330000 0.000000 2161.470000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.830000 0.000000 2156.970000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.330000 0.000000 2152.470000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830000 0.000000 2147.970000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.330000 0.000000 2143.470000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.830000 0.000000 2138.970000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.330000 0.000000 2134.470000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.830000 0.000000 2129.970000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.330000 0.000000 2125.470000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2120.830000 0.000000 2120.970000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2116.330000 0.000000 2116.470000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.830000 0.000000 2111.970000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.330000 0.000000 2107.470000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.830000 0.000000 2102.970000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.330000 0.000000 2098.470000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.730000 0.000000 2093.870000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.230000 0.000000 2089.370000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.730000 0.000000 2084.870000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.230000 0.000000 2080.370000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.730000 0.000000 2075.870000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.230000 0.000000 2071.370000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.730000 0.000000 2066.870000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.230000 0.000000 2062.370000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.730000 0.000000 2057.870000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.230000 0.000000 2053.370000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.730000 0.000000 2048.870000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.230000 0.000000 2044.370000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.730000 0.000000 2039.870000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.230000 0.000000 2035.370000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.730000 0.000000 2030.870000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.230000 0.000000 2026.370000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.730000 0.000000 2021.870000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.230000 0.000000 2017.370000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.730000 0.000000 2012.870000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.230000 0.000000 2008.370000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.730000 0.000000 2003.870000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.230000 0.000000 1999.370000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.730000 0.000000 1994.870000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.230000 0.000000 1990.370000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.730000 0.000000 1985.870000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.230000 0.000000 1981.370000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.730000 0.000000 1976.870000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.230000 0.000000 1972.370000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.730000 0.000000 1967.870000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.230000 0.000000 1963.370000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.730000 0.000000 1958.870000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.230000 0.000000 1954.370000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.730000 0.000000 1949.870000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.130000 0.000000 1945.270000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.630000 0.000000 1940.770000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.130000 0.000000 1936.270000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.630000 0.000000 1931.770000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.130000 0.000000 1927.270000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.630000 0.000000 1922.770000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.130000 0.000000 1918.270000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.630000 0.000000 1913.770000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.130000 0.000000 1909.270000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.630000 0.000000 1904.770000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.130000 0.000000 1900.270000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.630000 0.000000 1895.770000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.130000 0.000000 1891.270000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.630000 0.000000 1886.770000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.130000 0.000000 1882.270000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.630000 0.000000 1877.770000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.130000 0.000000 1873.270000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.630000 0.000000 1868.770000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.130000 0.000000 1864.270000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.630000 0.000000 1859.770000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.130000 0.000000 1855.270000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.630000 0.000000 1850.770000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.130000 0.000000 1846.270000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.630000 0.000000 1841.770000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.130000 0.000000 1837.270000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.630000 0.000000 1832.770000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.130000 0.000000 1828.270000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.630000 0.000000 1823.770000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.130000 0.000000 1819.270000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.630000 0.000000 1814.770000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.130000 0.000000 1810.270000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.630000 0.000000 1805.770000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.130000 0.000000 1801.270000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.530000 0.000000 1796.670000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.030000 0.000000 1792.170000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.530000 0.000000 1787.670000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.030000 0.000000 1783.170000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.530000 0.000000 1778.670000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.030000 0.000000 1774.170000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.530000 0.000000 1769.670000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.030000 0.000000 1765.170000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.530000 0.000000 1760.670000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.030000 0.000000 1756.170000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.530000 0.000000 1751.670000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.030000 0.000000 1747.170000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.530000 0.000000 1742.670000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.030000 0.000000 1738.170000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.530000 0.000000 1733.670000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.030000 0.000000 1729.170000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.530000 0.000000 1724.670000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.030000 0.000000 1720.170000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.530000 0.000000 1715.670000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.030000 0.000000 1711.170000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.530000 0.000000 1706.670000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.030000 0.000000 1702.170000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.530000 0.000000 1697.670000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.030000 0.000000 1693.170000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.530000 0.000000 1688.670000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.030000 0.000000 1684.170000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.530000 0.000000 1679.670000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.030000 0.000000 1675.170000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.530000 0.000000 1670.670000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.030000 0.000000 1666.170000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.530000 0.000000 1661.670000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.030000 0.000000 1657.170000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.530000 0.000000 1652.670000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.030000 0.000000 1648.170000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.430000 0.000000 1643.570000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.930000 0.000000 1639.070000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.430000 0.000000 1634.570000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.930000 0.000000 1630.070000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 71.660000 0.800000 71.960000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 179.415000 0.800000 179.715000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 287.250000 0.800000 287.550000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 430.955000 0.800000 431.255000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 574.655000 0.800000 574.955000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 718.355000 0.800000 718.655000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 862.135000 0.800000 862.435000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1005.755000 0.800000 1006.055000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1149.535000 0.800000 1149.835000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1293.240000 0.800000 1293.540000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1436.940000 0.800000 1437.240000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1580.720000 0.800000 1581.020000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1724.420000 0.800000 1724.720000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1868.120000 0.800000 1868.420000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.730000 2289.750000 126.870000 2290.240000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.530000 2289.750000 380.670000 2290.240000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.330000 2289.750000 634.470000 2290.240000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.030000 2289.750000 888.170000 2290.240000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.830000 2289.750000 1141.970000 2290.240000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.530000 2289.750000 1395.670000 2290.240000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.330000 2289.750000 1649.470000 2290.240000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.130000 2289.750000 1903.270000 2290.240000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.830000 2289.750000 2156.970000 2290.240000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1830.835000 2369.460000 1831.135000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1684.365000 2369.460000 1684.665000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1537.900000 2369.460000 1538.200000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1391.355000 2369.460000 1391.655000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1244.890000 2369.460000 1245.190000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1098.425000 2369.460000 1098.725000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 951.960000 2369.460000 952.260000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 805.415000 2369.460000 805.715000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 658.945000 2369.460000 659.245000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 549.060000 2369.460000 549.360000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 439.250000 2369.460000 439.550000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 329.360000 2369.460000 329.660000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 219.470000 2369.460000 219.770000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 109.580000 2369.460000 109.880000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1.590000 2369.460000 1.890000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2013.120000 0.800000 2013.420000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.470000 0.800000 143.770000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 251.305000 0.800000 251.605000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 395.010000 0.800000 395.310000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 538.710000 0.800000 539.010000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 682.490000 0.800000 682.790000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 826.110000 0.800000 826.410000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 969.890000 0.800000 970.190000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1113.590000 0.800000 1113.890000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1257.295000 0.800000 1257.595000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1400.995000 0.800000 1401.295000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1544.775000 0.800000 1545.075000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1688.475000 0.800000 1688.775000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1832.175000 0.800000 1832.475000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.330000 2289.750000 63.470000 2290.240000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.130000 2289.750000 317.270000 2290.240000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.830000 2289.750000 570.970000 2290.240000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.630000 2289.750000 824.770000 2290.240000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.330000 2289.750000 1078.470000 2290.240000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.130000 2289.750000 1332.270000 2290.240000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.930000 2289.750000 1586.070000 2290.240000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.630000 2289.750000 1839.770000 2290.240000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.430000 2289.750000 2093.570000 2290.240000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1867.410000 2369.460000 1867.710000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1720.945000 2369.460000 1721.245000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1574.480000 2369.460000 1574.780000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1428.010000 2369.460000 1428.310000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1281.465000 2369.460000 1281.765000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1135.000000 2369.460000 1135.300000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 988.535000 2369.460000 988.835000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 842.070000 2369.460000 842.370000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 695.525000 2369.460000 695.825000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 585.715000 2369.460000 586.015000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 475.905000 2369.460000 476.205000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 366.015000 2369.460000 366.315000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 256.125000 2369.460000 256.425000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 146.315000 2369.460000 146.615000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 36.425000 2369.460000 36.725000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2088.150000 0.800000 2088.450000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.525000 0.800000 107.825000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 215.360000 0.800000 215.660000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 359.065000 0.800000 359.365000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 502.765000 0.800000 503.065000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 646.545000 0.800000 646.845000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 790.245000 0.800000 790.545000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 933.945000 0.800000 934.245000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1077.725000 0.800000 1078.025000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1221.350000 0.800000 1221.650000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1365.130000 0.800000 1365.430000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1508.830000 0.800000 1509.130000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1652.530000 0.800000 1652.830000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1796.310000 0.800000 1796.610000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.330000 2289.750000 3.470000 2290.240000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.630000 2289.750000 253.770000 2290.240000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.430000 2289.750000 507.570000 2290.240000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.130000 2289.750000 761.270000 2290.240000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.930000 2289.750000 1015.070000 2290.240000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.730000 2289.750000 1268.870000 2290.240000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.430000 2289.750000 1522.570000 2290.240000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.230000 2289.750000 1776.370000 2290.240000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930000 2289.750000 2030.070000 2290.240000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1901.065000 2369.460000 1901.365000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1757.520000 2369.460000 1757.820000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1611.055000 2369.460000 1611.355000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1464.590000 2369.460000 1464.890000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1318.125000 2369.460000 1318.425000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1171.655000 2369.460000 1171.955000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1025.110000 2369.460000 1025.410000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 878.645000 2369.460000 878.945000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 732.180000 2369.460000 732.480000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 622.370000 2369.460000 622.670000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 512.480000 2369.460000 512.780000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 402.590000 2369.460000 402.890000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 292.780000 2369.460000 293.080000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 182.895000 2369.460000 183.195000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 73.005000 2369.460000 73.305000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.740000 0.000000 10.880000 0.485000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.140000 0.000000 6.280000 0.485000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.180000 0.595000 4.320000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2213.865000 1688.285000 2215.605000 2083.065000 ;
      LAYER met3 ;
        RECT 1738.545000 1688.285000 2215.605000 1690.025000 ;
      LAYER met3 ;
        RECT 1738.545000 2081.325000 2215.605000 2083.065000 ;
      LAYER met4 ;
        RECT 1738.545000 1688.285000 1740.285000 2083.065000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2213.865000 1222.785000 2215.605000 1617.565000 ;
      LAYER met3 ;
        RECT 1738.545000 1222.785000 2215.605000 1224.525000 ;
      LAYER met3 ;
        RECT 1738.545000 1615.825000 2215.605000 1617.565000 ;
      LAYER met4 ;
        RECT 1738.545000 1222.785000 1740.285000 1617.565000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2213.865000 757.285000 2215.605000 1152.065000 ;
      LAYER met3 ;
        RECT 1738.545000 757.285000 2215.605000 759.025000 ;
      LAYER met3 ;
        RECT 1738.545000 1150.325000 2215.605000 1152.065000 ;
      LAYER met4 ;
        RECT 1738.545000 757.285000 1740.285000 1152.065000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2213.865000 291.785000 2215.605000 686.565000 ;
      LAYER met3 ;
        RECT 1738.545000 291.785000 2215.605000 293.525000 ;
      LAYER met3 ;
        RECT 1738.545000 684.825000 2215.605000 686.565000 ;
      LAYER met4 ;
        RECT 1738.545000 291.785000 1740.285000 686.565000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 627.050000 1695.370000 628.790000 2090.150000 ;
      LAYER met3 ;
        RECT 151.730000 1695.370000 628.790000 1697.110000 ;
      LAYER met3 ;
        RECT 151.730000 2088.410000 628.790000 2090.150000 ;
      LAYER met4 ;
        RECT 151.730000 1695.370000 153.470000 2090.150000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 627.050000 1229.870000 628.790000 1624.650000 ;
      LAYER met3 ;
        RECT 151.730000 1229.870000 628.790000 1231.610000 ;
      LAYER met3 ;
        RECT 151.730000 1622.910000 628.790000 1624.650000 ;
      LAYER met4 ;
        RECT 151.730000 1229.870000 153.470000 1624.650000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 627.050000 764.370000 628.790000 1159.150000 ;
      LAYER met3 ;
        RECT 151.730000 764.370000 628.790000 766.110000 ;
      LAYER met3 ;
        RECT 151.730000 1157.410000 628.790000 1159.150000 ;
      LAYER met4 ;
        RECT 151.730000 764.370000 153.470000 1159.150000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 627.050000 298.870000 628.790000 693.650000 ;
      LAYER met3 ;
        RECT 151.730000 298.870000 628.790000 300.610000 ;
      LAYER met3 ;
        RECT 151.730000 691.910000 628.790000 693.650000 ;
      LAYER met4 ;
        RECT 151.730000 298.870000 153.470000 693.650000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1741.945000 2077.925000 2212.205000 2079.665000 ;
      LAYER met3 ;
        RECT 1741.945000 1691.685000 2212.205000 1693.425000 ;
      LAYER met4 ;
        RECT 1741.945000 1691.685000 1743.685000 2079.665000 ;
      LAYER met4 ;
        RECT 2210.465000 1691.685000 2212.205000 2079.665000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1741.945000 1612.425000 2212.205000 1614.165000 ;
      LAYER met3 ;
        RECT 1741.945000 1226.185000 2212.205000 1227.925000 ;
      LAYER met4 ;
        RECT 1741.945000 1226.185000 1743.685000 1614.165000 ;
      LAYER met4 ;
        RECT 2210.465000 1226.185000 2212.205000 1614.165000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1741.945000 1146.925000 2212.205000 1148.665000 ;
      LAYER met3 ;
        RECT 1741.945000 760.685000 2212.205000 762.425000 ;
      LAYER met4 ;
        RECT 1741.945000 760.685000 1743.685000 1148.665000 ;
      LAYER met4 ;
        RECT 2210.465000 760.685000 2212.205000 1148.665000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1741.945000 681.425000 2212.205000 683.165000 ;
      LAYER met3 ;
        RECT 1741.945000 295.185000 2212.205000 296.925000 ;
      LAYER met4 ;
        RECT 1741.945000 295.185000 1743.685000 683.165000 ;
      LAYER met4 ;
        RECT 2210.465000 295.185000 2212.205000 683.165000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 155.130000 2085.010000 625.390000 2086.750000 ;
      LAYER met3 ;
        RECT 155.130000 1698.770000 625.390000 1700.510000 ;
      LAYER met4 ;
        RECT 155.130000 1698.770000 156.870000 2086.750000 ;
      LAYER met4 ;
        RECT 623.650000 1698.770000 625.390000 2086.750000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 155.130000 1619.510000 625.390000 1621.250000 ;
      LAYER met3 ;
        RECT 155.130000 1233.270000 625.390000 1235.010000 ;
      LAYER met4 ;
        RECT 155.130000 1233.270000 156.870000 1621.250000 ;
      LAYER met4 ;
        RECT 623.650000 1233.270000 625.390000 1621.250000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 155.130000 1154.010000 625.390000 1155.750000 ;
      LAYER met3 ;
        RECT 155.130000 767.770000 625.390000 769.510000 ;
      LAYER met4 ;
        RECT 155.130000 767.770000 156.870000 1155.750000 ;
      LAYER met4 ;
        RECT 623.650000 767.770000 625.390000 1155.750000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 155.130000 688.510000 625.390000 690.250000 ;
      LAYER met3 ;
        RECT 155.130000 302.270000 625.390000 304.010000 ;
      LAYER met4 ;
        RECT 155.130000 302.270000 156.870000 690.250000 ;
      LAYER met4 ;
        RECT 623.650000 302.270000 625.390000 690.250000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2369.460000 2290.240000 ;
    LAYER met1 ;
      RECT 0.000000 4.460000 2369.460000 2290.240000 ;
      RECT 0.735000 4.040000 2369.460000 4.460000 ;
      RECT 0.000000 0.000000 2369.460000 4.040000 ;
    LAYER met2 ;
      RECT 2157.110000 2289.610000 2369.460000 2290.240000 ;
      RECT 2093.710000 2289.610000 2156.690000 2290.240000 ;
      RECT 2030.210000 2289.610000 2093.290000 2290.240000 ;
      RECT 1903.410000 2289.610000 2029.790000 2290.240000 ;
      RECT 1839.910000 2289.610000 1902.990000 2290.240000 ;
      RECT 1776.510000 2289.610000 1839.490000 2290.240000 ;
      RECT 1649.610000 2289.610000 1776.090000 2290.240000 ;
      RECT 1586.210000 2289.610000 1649.190000 2290.240000 ;
      RECT 1522.710000 2289.610000 1585.790000 2290.240000 ;
      RECT 1395.810000 2289.610000 1522.290000 2290.240000 ;
      RECT 1332.410000 2289.610000 1395.390000 2290.240000 ;
      RECT 1269.010000 2289.610000 1331.990000 2290.240000 ;
      RECT 1142.110000 2289.610000 1268.590000 2290.240000 ;
      RECT 1078.610000 2289.610000 1141.690000 2290.240000 ;
      RECT 1015.210000 2289.610000 1078.190000 2290.240000 ;
      RECT 888.310000 2289.610000 1014.790000 2290.240000 ;
      RECT 824.910000 2289.610000 887.890000 2290.240000 ;
      RECT 761.410000 2289.610000 824.490000 2290.240000 ;
      RECT 634.610000 2289.610000 760.990000 2290.240000 ;
      RECT 571.110000 2289.610000 634.190000 2290.240000 ;
      RECT 507.710000 2289.610000 570.690000 2290.240000 ;
      RECT 380.810000 2289.610000 507.290000 2290.240000 ;
      RECT 317.410000 2289.610000 380.390000 2290.240000 ;
      RECT 253.910000 2289.610000 316.990000 2290.240000 ;
      RECT 127.010000 2289.610000 253.490000 2290.240000 ;
      RECT 63.610000 2289.610000 126.590000 2290.240000 ;
      RECT 3.610000 2289.610000 63.190000 2290.240000 ;
      RECT 0.000000 2289.610000 3.190000 2290.240000 ;
      RECT 0.000000 0.630000 2369.460000 2289.610000 ;
      RECT 9.210000 0.625000 13.290000 0.630000 ;
      RECT 4.710000 0.625000 8.790000 0.630000 ;
      RECT 2202.110000 0.000000 2369.460000 0.630000 ;
      RECT 2197.610000 0.000000 2201.690000 0.630000 ;
      RECT 2193.110000 0.000000 2197.190000 0.630000 ;
      RECT 2188.610000 0.000000 2192.690000 0.630000 ;
      RECT 2184.110000 0.000000 2188.190000 0.630000 ;
      RECT 2179.610000 0.000000 2183.690000 0.630000 ;
      RECT 2175.110000 0.000000 2179.190000 0.630000 ;
      RECT 2170.610000 0.000000 2174.690000 0.630000 ;
      RECT 2166.110000 0.000000 2170.190000 0.630000 ;
      RECT 2161.610000 0.000000 2165.690000 0.630000 ;
      RECT 2157.110000 0.000000 2161.190000 0.630000 ;
      RECT 2152.610000 0.000000 2156.690000 0.630000 ;
      RECT 2148.110000 0.000000 2152.190000 0.630000 ;
      RECT 2143.610000 0.000000 2147.690000 0.630000 ;
      RECT 2139.110000 0.000000 2143.190000 0.630000 ;
      RECT 2134.610000 0.000000 2138.690000 0.630000 ;
      RECT 2130.110000 0.000000 2134.190000 0.630000 ;
      RECT 2125.610000 0.000000 2129.690000 0.630000 ;
      RECT 2121.110000 0.000000 2125.190000 0.630000 ;
      RECT 2116.610000 0.000000 2120.690000 0.630000 ;
      RECT 2112.110000 0.000000 2116.190000 0.630000 ;
      RECT 2107.610000 0.000000 2111.690000 0.630000 ;
      RECT 2103.110000 0.000000 2107.190000 0.630000 ;
      RECT 2098.610000 0.000000 2102.690000 0.630000 ;
      RECT 2094.010000 0.000000 2098.190000 0.630000 ;
      RECT 2089.510000 0.000000 2093.590000 0.630000 ;
      RECT 2085.010000 0.000000 2089.090000 0.630000 ;
      RECT 2080.510000 0.000000 2084.590000 0.630000 ;
      RECT 2076.010000 0.000000 2080.090000 0.630000 ;
      RECT 2071.510000 0.000000 2075.590000 0.630000 ;
      RECT 2067.010000 0.000000 2071.090000 0.630000 ;
      RECT 2062.510000 0.000000 2066.590000 0.630000 ;
      RECT 2058.010000 0.000000 2062.090000 0.630000 ;
      RECT 2053.510000 0.000000 2057.590000 0.630000 ;
      RECT 2049.010000 0.000000 2053.090000 0.630000 ;
      RECT 2044.510000 0.000000 2048.590000 0.630000 ;
      RECT 2040.010000 0.000000 2044.090000 0.630000 ;
      RECT 2035.510000 0.000000 2039.590000 0.630000 ;
      RECT 2031.010000 0.000000 2035.090000 0.630000 ;
      RECT 2026.510000 0.000000 2030.590000 0.630000 ;
      RECT 2022.010000 0.000000 2026.090000 0.630000 ;
      RECT 2017.510000 0.000000 2021.590000 0.630000 ;
      RECT 2013.010000 0.000000 2017.090000 0.630000 ;
      RECT 2008.510000 0.000000 2012.590000 0.630000 ;
      RECT 2004.010000 0.000000 2008.090000 0.630000 ;
      RECT 1999.510000 0.000000 2003.590000 0.630000 ;
      RECT 1995.010000 0.000000 1999.090000 0.630000 ;
      RECT 1990.510000 0.000000 1994.590000 0.630000 ;
      RECT 1986.010000 0.000000 1990.090000 0.630000 ;
      RECT 1981.510000 0.000000 1985.590000 0.630000 ;
      RECT 1977.010000 0.000000 1981.090000 0.630000 ;
      RECT 1972.510000 0.000000 1976.590000 0.630000 ;
      RECT 1968.010000 0.000000 1972.090000 0.630000 ;
      RECT 1963.510000 0.000000 1967.590000 0.630000 ;
      RECT 1959.010000 0.000000 1963.090000 0.630000 ;
      RECT 1954.510000 0.000000 1958.590000 0.630000 ;
      RECT 1950.010000 0.000000 1954.090000 0.630000 ;
      RECT 1945.410000 0.000000 1949.590000 0.630000 ;
      RECT 1940.910000 0.000000 1944.990000 0.630000 ;
      RECT 1936.410000 0.000000 1940.490000 0.630000 ;
      RECT 1931.910000 0.000000 1935.990000 0.630000 ;
      RECT 1927.410000 0.000000 1931.490000 0.630000 ;
      RECT 1922.910000 0.000000 1926.990000 0.630000 ;
      RECT 1918.410000 0.000000 1922.490000 0.630000 ;
      RECT 1913.910000 0.000000 1917.990000 0.630000 ;
      RECT 1909.410000 0.000000 1913.490000 0.630000 ;
      RECT 1904.910000 0.000000 1908.990000 0.630000 ;
      RECT 1900.410000 0.000000 1904.490000 0.630000 ;
      RECT 1895.910000 0.000000 1899.990000 0.630000 ;
      RECT 1891.410000 0.000000 1895.490000 0.630000 ;
      RECT 1886.910000 0.000000 1890.990000 0.630000 ;
      RECT 1882.410000 0.000000 1886.490000 0.630000 ;
      RECT 1877.910000 0.000000 1881.990000 0.630000 ;
      RECT 1873.410000 0.000000 1877.490000 0.630000 ;
      RECT 1868.910000 0.000000 1872.990000 0.630000 ;
      RECT 1864.410000 0.000000 1868.490000 0.630000 ;
      RECT 1859.910000 0.000000 1863.990000 0.630000 ;
      RECT 1855.410000 0.000000 1859.490000 0.630000 ;
      RECT 1850.910000 0.000000 1854.990000 0.630000 ;
      RECT 1846.410000 0.000000 1850.490000 0.630000 ;
      RECT 1841.910000 0.000000 1845.990000 0.630000 ;
      RECT 1837.410000 0.000000 1841.490000 0.630000 ;
      RECT 1832.910000 0.000000 1836.990000 0.630000 ;
      RECT 1828.410000 0.000000 1832.490000 0.630000 ;
      RECT 1823.910000 0.000000 1827.990000 0.630000 ;
      RECT 1819.410000 0.000000 1823.490000 0.630000 ;
      RECT 1814.910000 0.000000 1818.990000 0.630000 ;
      RECT 1810.410000 0.000000 1814.490000 0.630000 ;
      RECT 1805.910000 0.000000 1809.990000 0.630000 ;
      RECT 1801.410000 0.000000 1805.490000 0.630000 ;
      RECT 1796.810000 0.000000 1800.990000 0.630000 ;
      RECT 1792.310000 0.000000 1796.390000 0.630000 ;
      RECT 1787.810000 0.000000 1791.890000 0.630000 ;
      RECT 1783.310000 0.000000 1787.390000 0.630000 ;
      RECT 1778.810000 0.000000 1782.890000 0.630000 ;
      RECT 1774.310000 0.000000 1778.390000 0.630000 ;
      RECT 1769.810000 0.000000 1773.890000 0.630000 ;
      RECT 1765.310000 0.000000 1769.390000 0.630000 ;
      RECT 1760.810000 0.000000 1764.890000 0.630000 ;
      RECT 1756.310000 0.000000 1760.390000 0.630000 ;
      RECT 1751.810000 0.000000 1755.890000 0.630000 ;
      RECT 1747.310000 0.000000 1751.390000 0.630000 ;
      RECT 1742.810000 0.000000 1746.890000 0.630000 ;
      RECT 1738.310000 0.000000 1742.390000 0.630000 ;
      RECT 1733.810000 0.000000 1737.890000 0.630000 ;
      RECT 1729.310000 0.000000 1733.390000 0.630000 ;
      RECT 1724.810000 0.000000 1728.890000 0.630000 ;
      RECT 1720.310000 0.000000 1724.390000 0.630000 ;
      RECT 1715.810000 0.000000 1719.890000 0.630000 ;
      RECT 1711.310000 0.000000 1715.390000 0.630000 ;
      RECT 1706.810000 0.000000 1710.890000 0.630000 ;
      RECT 1702.310000 0.000000 1706.390000 0.630000 ;
      RECT 1697.810000 0.000000 1701.890000 0.630000 ;
      RECT 1693.310000 0.000000 1697.390000 0.630000 ;
      RECT 1688.810000 0.000000 1692.890000 0.630000 ;
      RECT 1684.310000 0.000000 1688.390000 0.630000 ;
      RECT 1679.810000 0.000000 1683.890000 0.630000 ;
      RECT 1675.310000 0.000000 1679.390000 0.630000 ;
      RECT 1670.810000 0.000000 1674.890000 0.630000 ;
      RECT 1666.310000 0.000000 1670.390000 0.630000 ;
      RECT 1661.810000 0.000000 1665.890000 0.630000 ;
      RECT 1657.310000 0.000000 1661.390000 0.630000 ;
      RECT 1652.810000 0.000000 1656.890000 0.630000 ;
      RECT 1648.310000 0.000000 1652.390000 0.630000 ;
      RECT 1643.710000 0.000000 1647.890000 0.630000 ;
      RECT 1639.210000 0.000000 1643.290000 0.630000 ;
      RECT 1634.710000 0.000000 1638.790000 0.630000 ;
      RECT 1630.210000 0.000000 1634.290000 0.630000 ;
      RECT 1625.710000 0.000000 1629.790000 0.630000 ;
      RECT 1621.210000 0.000000 1625.290000 0.630000 ;
      RECT 1616.710000 0.000000 1620.790000 0.630000 ;
      RECT 1612.210000 0.000000 1616.290000 0.630000 ;
      RECT 1607.710000 0.000000 1611.790000 0.630000 ;
      RECT 1603.210000 0.000000 1607.290000 0.630000 ;
      RECT 1598.710000 0.000000 1602.790000 0.630000 ;
      RECT 1594.210000 0.000000 1598.290000 0.630000 ;
      RECT 1589.710000 0.000000 1593.790000 0.630000 ;
      RECT 1585.210000 0.000000 1589.290000 0.630000 ;
      RECT 1580.710000 0.000000 1584.790000 0.630000 ;
      RECT 1576.210000 0.000000 1580.290000 0.630000 ;
      RECT 1571.710000 0.000000 1575.790000 0.630000 ;
      RECT 1567.210000 0.000000 1571.290000 0.630000 ;
      RECT 1562.710000 0.000000 1566.790000 0.630000 ;
      RECT 1558.210000 0.000000 1562.290000 0.630000 ;
      RECT 1553.710000 0.000000 1557.790000 0.630000 ;
      RECT 1549.210000 0.000000 1553.290000 0.630000 ;
      RECT 1544.710000 0.000000 1548.790000 0.630000 ;
      RECT 1540.210000 0.000000 1544.290000 0.630000 ;
      RECT 1535.710000 0.000000 1539.790000 0.630000 ;
      RECT 1531.210000 0.000000 1535.290000 0.630000 ;
      RECT 1526.710000 0.000000 1530.790000 0.630000 ;
      RECT 1522.210000 0.000000 1526.290000 0.630000 ;
      RECT 1517.710000 0.000000 1521.790000 0.630000 ;
      RECT 1513.210000 0.000000 1517.290000 0.630000 ;
      RECT 1508.710000 0.000000 1512.790000 0.630000 ;
      RECT 1504.210000 0.000000 1508.290000 0.630000 ;
      RECT 1499.710000 0.000000 1503.790000 0.630000 ;
      RECT 1495.110000 0.000000 1499.290000 0.630000 ;
      RECT 1490.610000 0.000000 1494.690000 0.630000 ;
      RECT 1486.110000 0.000000 1490.190000 0.630000 ;
      RECT 1481.610000 0.000000 1485.690000 0.630000 ;
      RECT 1477.110000 0.000000 1481.190000 0.630000 ;
      RECT 1472.610000 0.000000 1476.690000 0.630000 ;
      RECT 1468.110000 0.000000 1472.190000 0.630000 ;
      RECT 1463.610000 0.000000 1467.690000 0.630000 ;
      RECT 1459.110000 0.000000 1463.190000 0.630000 ;
      RECT 1454.610000 0.000000 1458.690000 0.630000 ;
      RECT 1450.110000 0.000000 1454.190000 0.630000 ;
      RECT 1445.610000 0.000000 1449.690000 0.630000 ;
      RECT 1441.110000 0.000000 1445.190000 0.630000 ;
      RECT 1436.610000 0.000000 1440.690000 0.630000 ;
      RECT 1432.110000 0.000000 1436.190000 0.630000 ;
      RECT 1427.610000 0.000000 1431.690000 0.630000 ;
      RECT 1423.110000 0.000000 1427.190000 0.630000 ;
      RECT 1418.610000 0.000000 1422.690000 0.630000 ;
      RECT 1414.110000 0.000000 1418.190000 0.630000 ;
      RECT 1409.610000 0.000000 1413.690000 0.630000 ;
      RECT 1405.110000 0.000000 1409.190000 0.630000 ;
      RECT 1400.610000 0.000000 1404.690000 0.630000 ;
      RECT 1396.110000 0.000000 1400.190000 0.630000 ;
      RECT 1391.610000 0.000000 1395.690000 0.630000 ;
      RECT 1387.110000 0.000000 1391.190000 0.630000 ;
      RECT 1382.610000 0.000000 1386.690000 0.630000 ;
      RECT 1378.110000 0.000000 1382.190000 0.630000 ;
      RECT 1373.610000 0.000000 1377.690000 0.630000 ;
      RECT 1369.110000 0.000000 1373.190000 0.630000 ;
      RECT 1364.610000 0.000000 1368.690000 0.630000 ;
      RECT 1360.110000 0.000000 1364.190000 0.630000 ;
      RECT 1355.610000 0.000000 1359.690000 0.630000 ;
      RECT 1351.110000 0.000000 1355.190000 0.630000 ;
      RECT 1346.510000 0.000000 1350.690000 0.630000 ;
      RECT 1342.010000 0.000000 1346.090000 0.630000 ;
      RECT 1337.510000 0.000000 1341.590000 0.630000 ;
      RECT 1333.010000 0.000000 1337.090000 0.630000 ;
      RECT 1328.510000 0.000000 1332.590000 0.630000 ;
      RECT 1324.010000 0.000000 1328.090000 0.630000 ;
      RECT 1319.510000 0.000000 1323.590000 0.630000 ;
      RECT 1315.010000 0.000000 1319.090000 0.630000 ;
      RECT 1310.510000 0.000000 1314.590000 0.630000 ;
      RECT 1306.010000 0.000000 1310.090000 0.630000 ;
      RECT 1301.510000 0.000000 1305.590000 0.630000 ;
      RECT 1297.010000 0.000000 1301.090000 0.630000 ;
      RECT 1292.510000 0.000000 1296.590000 0.630000 ;
      RECT 1288.010000 0.000000 1292.090000 0.630000 ;
      RECT 1283.510000 0.000000 1287.590000 0.630000 ;
      RECT 1279.010000 0.000000 1283.090000 0.630000 ;
      RECT 1274.510000 0.000000 1278.590000 0.630000 ;
      RECT 1270.010000 0.000000 1274.090000 0.630000 ;
      RECT 1265.510000 0.000000 1269.590000 0.630000 ;
      RECT 1261.010000 0.000000 1265.090000 0.630000 ;
      RECT 1256.510000 0.000000 1260.590000 0.630000 ;
      RECT 1252.010000 0.000000 1256.090000 0.630000 ;
      RECT 1247.510000 0.000000 1251.590000 0.630000 ;
      RECT 1243.010000 0.000000 1247.090000 0.630000 ;
      RECT 1238.510000 0.000000 1242.590000 0.630000 ;
      RECT 1234.010000 0.000000 1238.090000 0.630000 ;
      RECT 1229.510000 0.000000 1233.590000 0.630000 ;
      RECT 1225.010000 0.000000 1229.090000 0.630000 ;
      RECT 1220.510000 0.000000 1224.590000 0.630000 ;
      RECT 1216.010000 0.000000 1220.090000 0.630000 ;
      RECT 1211.510000 0.000000 1215.590000 0.630000 ;
      RECT 1207.010000 0.000000 1211.090000 0.630000 ;
      RECT 1202.510000 0.000000 1206.590000 0.630000 ;
      RECT 1198.010000 0.000000 1202.090000 0.630000 ;
      RECT 1193.410000 0.000000 1197.590000 0.630000 ;
      RECT 1188.910000 0.000000 1192.990000 0.630000 ;
      RECT 1184.410000 0.000000 1188.490000 0.630000 ;
      RECT 1179.910000 0.000000 1183.990000 0.630000 ;
      RECT 1175.410000 0.000000 1179.490000 0.630000 ;
      RECT 1170.910000 0.000000 1174.990000 0.630000 ;
      RECT 1166.410000 0.000000 1170.490000 0.630000 ;
      RECT 1161.910000 0.000000 1165.990000 0.630000 ;
      RECT 1157.410000 0.000000 1161.490000 0.630000 ;
      RECT 1152.910000 0.000000 1156.990000 0.630000 ;
      RECT 1148.410000 0.000000 1152.490000 0.630000 ;
      RECT 1143.910000 0.000000 1147.990000 0.630000 ;
      RECT 1139.410000 0.000000 1143.490000 0.630000 ;
      RECT 1134.910000 0.000000 1138.990000 0.630000 ;
      RECT 1130.410000 0.000000 1134.490000 0.630000 ;
      RECT 1125.910000 0.000000 1129.990000 0.630000 ;
      RECT 1121.410000 0.000000 1125.490000 0.630000 ;
      RECT 1116.910000 0.000000 1120.990000 0.630000 ;
      RECT 1112.410000 0.000000 1116.490000 0.630000 ;
      RECT 1107.910000 0.000000 1111.990000 0.630000 ;
      RECT 1103.410000 0.000000 1107.490000 0.630000 ;
      RECT 1098.910000 0.000000 1102.990000 0.630000 ;
      RECT 1094.410000 0.000000 1098.490000 0.630000 ;
      RECT 1089.910000 0.000000 1093.990000 0.630000 ;
      RECT 1085.410000 0.000000 1089.490000 0.630000 ;
      RECT 1080.910000 0.000000 1084.990000 0.630000 ;
      RECT 1076.410000 0.000000 1080.490000 0.630000 ;
      RECT 1071.910000 0.000000 1075.990000 0.630000 ;
      RECT 1067.410000 0.000000 1071.490000 0.630000 ;
      RECT 1062.910000 0.000000 1066.990000 0.630000 ;
      RECT 1058.410000 0.000000 1062.490000 0.630000 ;
      RECT 1053.910000 0.000000 1057.990000 0.630000 ;
      RECT 1049.410000 0.000000 1053.490000 0.630000 ;
      RECT 1044.810000 0.000000 1048.990000 0.630000 ;
      RECT 1040.310000 0.000000 1044.390000 0.630000 ;
      RECT 1035.810000 0.000000 1039.890000 0.630000 ;
      RECT 1031.310000 0.000000 1035.390000 0.630000 ;
      RECT 1026.810000 0.000000 1030.890000 0.630000 ;
      RECT 1022.310000 0.000000 1026.390000 0.630000 ;
      RECT 1017.810000 0.000000 1021.890000 0.630000 ;
      RECT 1013.310000 0.000000 1017.390000 0.630000 ;
      RECT 1008.810000 0.000000 1012.890000 0.630000 ;
      RECT 1004.310000 0.000000 1008.390000 0.630000 ;
      RECT 999.810000 0.000000 1003.890000 0.630000 ;
      RECT 995.310000 0.000000 999.390000 0.630000 ;
      RECT 990.810000 0.000000 994.890000 0.630000 ;
      RECT 986.310000 0.000000 990.390000 0.630000 ;
      RECT 981.810000 0.000000 985.890000 0.630000 ;
      RECT 977.310000 0.000000 981.390000 0.630000 ;
      RECT 972.810000 0.000000 976.890000 0.630000 ;
      RECT 968.310000 0.000000 972.390000 0.630000 ;
      RECT 963.810000 0.000000 967.890000 0.630000 ;
      RECT 959.310000 0.000000 963.390000 0.630000 ;
      RECT 954.810000 0.000000 958.890000 0.630000 ;
      RECT 950.310000 0.000000 954.390000 0.630000 ;
      RECT 945.810000 0.000000 949.890000 0.630000 ;
      RECT 941.310000 0.000000 945.390000 0.630000 ;
      RECT 936.810000 0.000000 940.890000 0.630000 ;
      RECT 932.310000 0.000000 936.390000 0.630000 ;
      RECT 927.810000 0.000000 931.890000 0.630000 ;
      RECT 923.310000 0.000000 927.390000 0.630000 ;
      RECT 918.810000 0.000000 922.890000 0.630000 ;
      RECT 914.310000 0.000000 918.390000 0.630000 ;
      RECT 909.810000 0.000000 913.890000 0.630000 ;
      RECT 905.310000 0.000000 909.390000 0.630000 ;
      RECT 900.810000 0.000000 904.890000 0.630000 ;
      RECT 896.210000 0.000000 900.390000 0.630000 ;
      RECT 891.710000 0.000000 895.790000 0.630000 ;
      RECT 887.210000 0.000000 891.290000 0.630000 ;
      RECT 882.710000 0.000000 886.790000 0.630000 ;
      RECT 878.210000 0.000000 882.290000 0.630000 ;
      RECT 873.710000 0.000000 877.790000 0.630000 ;
      RECT 869.210000 0.000000 873.290000 0.630000 ;
      RECT 864.710000 0.000000 868.790000 0.630000 ;
      RECT 860.210000 0.000000 864.290000 0.630000 ;
      RECT 855.710000 0.000000 859.790000 0.630000 ;
      RECT 851.210000 0.000000 855.290000 0.630000 ;
      RECT 846.710000 0.000000 850.790000 0.630000 ;
      RECT 842.210000 0.000000 846.290000 0.630000 ;
      RECT 837.710000 0.000000 841.790000 0.630000 ;
      RECT 833.210000 0.000000 837.290000 0.630000 ;
      RECT 828.710000 0.000000 832.790000 0.630000 ;
      RECT 824.210000 0.000000 828.290000 0.630000 ;
      RECT 819.710000 0.000000 823.790000 0.630000 ;
      RECT 815.210000 0.000000 819.290000 0.630000 ;
      RECT 810.710000 0.000000 814.790000 0.630000 ;
      RECT 806.210000 0.000000 810.290000 0.630000 ;
      RECT 801.710000 0.000000 805.790000 0.630000 ;
      RECT 797.210000 0.000000 801.290000 0.630000 ;
      RECT 792.710000 0.000000 796.790000 0.630000 ;
      RECT 788.210000 0.000000 792.290000 0.630000 ;
      RECT 783.710000 0.000000 787.790000 0.630000 ;
      RECT 779.210000 0.000000 783.290000 0.630000 ;
      RECT 774.710000 0.000000 778.790000 0.630000 ;
      RECT 770.210000 0.000000 774.290000 0.630000 ;
      RECT 765.710000 0.000000 769.790000 0.630000 ;
      RECT 761.210000 0.000000 765.290000 0.630000 ;
      RECT 756.710000 0.000000 760.790000 0.630000 ;
      RECT 752.210000 0.000000 756.290000 0.630000 ;
      RECT 747.710000 0.000000 751.790000 0.630000 ;
      RECT 743.110000 0.000000 747.290000 0.630000 ;
      RECT 738.610000 0.000000 742.690000 0.630000 ;
      RECT 734.110000 0.000000 738.190000 0.630000 ;
      RECT 729.610000 0.000000 733.690000 0.630000 ;
      RECT 725.110000 0.000000 729.190000 0.630000 ;
      RECT 720.610000 0.000000 724.690000 0.630000 ;
      RECT 716.110000 0.000000 720.190000 0.630000 ;
      RECT 711.610000 0.000000 715.690000 0.630000 ;
      RECT 707.110000 0.000000 711.190000 0.630000 ;
      RECT 702.610000 0.000000 706.690000 0.630000 ;
      RECT 698.110000 0.000000 702.190000 0.630000 ;
      RECT 693.610000 0.000000 697.690000 0.630000 ;
      RECT 689.110000 0.000000 693.190000 0.630000 ;
      RECT 684.610000 0.000000 688.690000 0.630000 ;
      RECT 680.110000 0.000000 684.190000 0.630000 ;
      RECT 675.610000 0.000000 679.690000 0.630000 ;
      RECT 671.110000 0.000000 675.190000 0.630000 ;
      RECT 666.610000 0.000000 670.690000 0.630000 ;
      RECT 662.110000 0.000000 666.190000 0.630000 ;
      RECT 657.610000 0.000000 661.690000 0.630000 ;
      RECT 653.110000 0.000000 657.190000 0.630000 ;
      RECT 648.610000 0.000000 652.690000 0.630000 ;
      RECT 644.110000 0.000000 648.190000 0.630000 ;
      RECT 639.610000 0.000000 643.690000 0.630000 ;
      RECT 635.110000 0.000000 639.190000 0.630000 ;
      RECT 630.610000 0.000000 634.690000 0.630000 ;
      RECT 626.110000 0.000000 630.190000 0.630000 ;
      RECT 621.610000 0.000000 625.690000 0.630000 ;
      RECT 617.110000 0.000000 621.190000 0.630000 ;
      RECT 612.610000 0.000000 616.690000 0.630000 ;
      RECT 608.110000 0.000000 612.190000 0.630000 ;
      RECT 603.610000 0.000000 607.690000 0.630000 ;
      RECT 599.110000 0.000000 603.190000 0.630000 ;
      RECT 594.510000 0.000000 598.690000 0.630000 ;
      RECT 590.010000 0.000000 594.090000 0.630000 ;
      RECT 585.510000 0.000000 589.590000 0.630000 ;
      RECT 581.010000 0.000000 585.090000 0.630000 ;
      RECT 576.510000 0.000000 580.590000 0.630000 ;
      RECT 572.010000 0.000000 576.090000 0.630000 ;
      RECT 567.510000 0.000000 571.590000 0.630000 ;
      RECT 563.010000 0.000000 567.090000 0.630000 ;
      RECT 558.510000 0.000000 562.590000 0.630000 ;
      RECT 554.010000 0.000000 558.090000 0.630000 ;
      RECT 549.510000 0.000000 553.590000 0.630000 ;
      RECT 545.010000 0.000000 549.090000 0.630000 ;
      RECT 540.510000 0.000000 544.590000 0.630000 ;
      RECT 536.010000 0.000000 540.090000 0.630000 ;
      RECT 531.510000 0.000000 535.590000 0.630000 ;
      RECT 527.010000 0.000000 531.090000 0.630000 ;
      RECT 522.510000 0.000000 526.590000 0.630000 ;
      RECT 518.010000 0.000000 522.090000 0.630000 ;
      RECT 513.510000 0.000000 517.590000 0.630000 ;
      RECT 509.010000 0.000000 513.090000 0.630000 ;
      RECT 504.510000 0.000000 508.590000 0.630000 ;
      RECT 500.010000 0.000000 504.090000 0.630000 ;
      RECT 495.510000 0.000000 499.590000 0.630000 ;
      RECT 491.010000 0.000000 495.090000 0.630000 ;
      RECT 486.510000 0.000000 490.590000 0.630000 ;
      RECT 482.010000 0.000000 486.090000 0.630000 ;
      RECT 477.510000 0.000000 481.590000 0.630000 ;
      RECT 473.010000 0.000000 477.090000 0.630000 ;
      RECT 468.510000 0.000000 472.590000 0.630000 ;
      RECT 464.010000 0.000000 468.090000 0.630000 ;
      RECT 459.510000 0.000000 463.590000 0.630000 ;
      RECT 455.010000 0.000000 459.090000 0.630000 ;
      RECT 450.510000 0.000000 454.590000 0.630000 ;
      RECT 445.910000 0.000000 450.090000 0.630000 ;
      RECT 441.410000 0.000000 445.490000 0.630000 ;
      RECT 436.910000 0.000000 440.990000 0.630000 ;
      RECT 432.410000 0.000000 436.490000 0.630000 ;
      RECT 427.910000 0.000000 431.990000 0.630000 ;
      RECT 423.410000 0.000000 427.490000 0.630000 ;
      RECT 418.910000 0.000000 422.990000 0.630000 ;
      RECT 414.410000 0.000000 418.490000 0.630000 ;
      RECT 409.910000 0.000000 413.990000 0.630000 ;
      RECT 405.410000 0.000000 409.490000 0.630000 ;
      RECT 400.910000 0.000000 404.990000 0.630000 ;
      RECT 396.410000 0.000000 400.490000 0.630000 ;
      RECT 391.910000 0.000000 395.990000 0.630000 ;
      RECT 387.410000 0.000000 391.490000 0.630000 ;
      RECT 382.910000 0.000000 386.990000 0.630000 ;
      RECT 378.410000 0.000000 382.490000 0.630000 ;
      RECT 373.910000 0.000000 377.990000 0.630000 ;
      RECT 369.410000 0.000000 373.490000 0.630000 ;
      RECT 364.910000 0.000000 368.990000 0.630000 ;
      RECT 360.410000 0.000000 364.490000 0.630000 ;
      RECT 355.910000 0.000000 359.990000 0.630000 ;
      RECT 351.410000 0.000000 355.490000 0.630000 ;
      RECT 346.910000 0.000000 350.990000 0.630000 ;
      RECT 342.410000 0.000000 346.490000 0.630000 ;
      RECT 337.910000 0.000000 341.990000 0.630000 ;
      RECT 333.410000 0.000000 337.490000 0.630000 ;
      RECT 328.910000 0.000000 332.990000 0.630000 ;
      RECT 324.410000 0.000000 328.490000 0.630000 ;
      RECT 319.910000 0.000000 323.990000 0.630000 ;
      RECT 315.410000 0.000000 319.490000 0.630000 ;
      RECT 310.910000 0.000000 314.990000 0.630000 ;
      RECT 306.410000 0.000000 310.490000 0.630000 ;
      RECT 301.910000 0.000000 305.990000 0.630000 ;
      RECT 297.410000 0.000000 301.490000 0.630000 ;
      RECT 292.810000 0.000000 296.990000 0.630000 ;
      RECT 288.310000 0.000000 292.390000 0.630000 ;
      RECT 283.810000 0.000000 287.890000 0.630000 ;
      RECT 279.310000 0.000000 283.390000 0.630000 ;
      RECT 274.810000 0.000000 278.890000 0.630000 ;
      RECT 270.310000 0.000000 274.390000 0.630000 ;
      RECT 265.810000 0.000000 269.890000 0.630000 ;
      RECT 261.310000 0.000000 265.390000 0.630000 ;
      RECT 256.810000 0.000000 260.890000 0.630000 ;
      RECT 252.310000 0.000000 256.390000 0.630000 ;
      RECT 247.810000 0.000000 251.890000 0.630000 ;
      RECT 243.310000 0.000000 247.390000 0.630000 ;
      RECT 238.810000 0.000000 242.890000 0.630000 ;
      RECT 234.310000 0.000000 238.390000 0.630000 ;
      RECT 229.810000 0.000000 233.890000 0.630000 ;
      RECT 225.310000 0.000000 229.390000 0.630000 ;
      RECT 220.810000 0.000000 224.890000 0.630000 ;
      RECT 216.310000 0.000000 220.390000 0.630000 ;
      RECT 211.810000 0.000000 215.890000 0.630000 ;
      RECT 207.310000 0.000000 211.390000 0.630000 ;
      RECT 202.810000 0.000000 206.890000 0.630000 ;
      RECT 198.310000 0.000000 202.390000 0.630000 ;
      RECT 193.810000 0.000000 197.890000 0.630000 ;
      RECT 189.310000 0.000000 193.390000 0.630000 ;
      RECT 184.810000 0.000000 188.890000 0.630000 ;
      RECT 180.310000 0.000000 184.390000 0.630000 ;
      RECT 175.810000 0.000000 179.890000 0.630000 ;
      RECT 171.310000 0.000000 175.390000 0.630000 ;
      RECT 166.810000 0.000000 170.890000 0.630000 ;
      RECT 162.310000 0.000000 166.390000 0.630000 ;
      RECT 157.810000 0.000000 161.890000 0.630000 ;
      RECT 153.310000 0.000000 157.390000 0.630000 ;
      RECT 148.810000 0.000000 152.890000 0.630000 ;
      RECT 144.210000 0.000000 148.390000 0.630000 ;
      RECT 139.710000 0.000000 143.790000 0.630000 ;
      RECT 135.210000 0.000000 139.290000 0.630000 ;
      RECT 130.710000 0.000000 134.790000 0.630000 ;
      RECT 126.210000 0.000000 130.290000 0.630000 ;
      RECT 121.710000 0.000000 125.790000 0.630000 ;
      RECT 117.210000 0.000000 121.290000 0.630000 ;
      RECT 112.710000 0.000000 116.790000 0.630000 ;
      RECT 108.210000 0.000000 112.290000 0.630000 ;
      RECT 103.710000 0.000000 107.790000 0.630000 ;
      RECT 99.210000 0.000000 103.290000 0.630000 ;
      RECT 94.710000 0.000000 98.790000 0.630000 ;
      RECT 90.210000 0.000000 94.290000 0.630000 ;
      RECT 85.710000 0.000000 89.790000 0.630000 ;
      RECT 81.210000 0.000000 85.290000 0.630000 ;
      RECT 76.710000 0.000000 80.790000 0.630000 ;
      RECT 72.210000 0.000000 76.290000 0.630000 ;
      RECT 67.710000 0.000000 71.790000 0.630000 ;
      RECT 63.210000 0.000000 67.290000 0.630000 ;
      RECT 58.710000 0.000000 62.790000 0.630000 ;
      RECT 54.210000 0.000000 58.290000 0.630000 ;
      RECT 49.710000 0.000000 53.790000 0.630000 ;
      RECT 45.210000 0.000000 49.290000 0.630000 ;
      RECT 40.710000 0.000000 44.790000 0.630000 ;
      RECT 36.210000 0.000000 40.290000 0.630000 ;
      RECT 31.710000 0.000000 35.790000 0.630000 ;
      RECT 27.210000 0.000000 31.290000 0.630000 ;
      RECT 22.710000 0.000000 26.790000 0.630000 ;
      RECT 18.210000 0.000000 22.290000 0.630000 ;
      RECT 13.710000 0.000000 17.790000 0.630000 ;
      RECT 11.020000 0.000000 13.290000 0.625000 ;
      RECT 9.210000 0.000000 10.600000 0.625000 ;
      RECT 6.420000 0.000000 8.790000 0.625000 ;
      RECT 4.710000 0.000000 6.000000 0.625000 ;
      RECT 1.810000 0.000000 4.290000 0.630000 ;
      RECT 0.000000 0.000000 1.390000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 2088.750000 2369.460000 2290.240000 ;
      RECT 1.100000 2087.850000 2369.460000 2088.750000 ;
      RECT 0.000000 2013.720000 2369.460000 2087.850000 ;
      RECT 1.100000 2012.820000 2369.460000 2013.720000 ;
      RECT 0.000000 1901.665000 2369.460000 2012.820000 ;
      RECT 0.000000 1900.765000 2368.360000 1901.665000 ;
      RECT 0.000000 1868.720000 2369.460000 1900.765000 ;
      RECT 1.100000 1868.010000 2369.460000 1868.720000 ;
      RECT 1.100000 1867.820000 2368.360000 1868.010000 ;
      RECT 0.000000 1867.110000 2368.360000 1867.820000 ;
      RECT 0.000000 1832.775000 2369.460000 1867.110000 ;
      RECT 1.100000 1831.875000 2369.460000 1832.775000 ;
      RECT 0.000000 1831.435000 2369.460000 1831.875000 ;
      RECT 0.000000 1830.535000 2368.360000 1831.435000 ;
      RECT 0.000000 1796.910000 2369.460000 1830.535000 ;
      RECT 1.100000 1796.010000 2369.460000 1796.910000 ;
      RECT 0.000000 1758.120000 2369.460000 1796.010000 ;
      RECT 0.000000 1757.220000 2368.360000 1758.120000 ;
      RECT 0.000000 1725.020000 2369.460000 1757.220000 ;
      RECT 1.100000 1724.120000 2369.460000 1725.020000 ;
      RECT 0.000000 1721.545000 2369.460000 1724.120000 ;
      RECT 0.000000 1720.645000 2368.360000 1721.545000 ;
      RECT 0.000000 1689.075000 2369.460000 1720.645000 ;
      RECT 1.100000 1688.175000 2369.460000 1689.075000 ;
      RECT 0.000000 1684.965000 2369.460000 1688.175000 ;
      RECT 0.000000 1684.065000 2368.360000 1684.965000 ;
      RECT 0.000000 1653.130000 2369.460000 1684.065000 ;
      RECT 1.100000 1652.230000 2369.460000 1653.130000 ;
      RECT 0.000000 1611.655000 2369.460000 1652.230000 ;
      RECT 0.000000 1610.755000 2368.360000 1611.655000 ;
      RECT 0.000000 1581.320000 2369.460000 1610.755000 ;
      RECT 1.100000 1580.420000 2369.460000 1581.320000 ;
      RECT 0.000000 1575.080000 2369.460000 1580.420000 ;
      RECT 0.000000 1574.180000 2368.360000 1575.080000 ;
      RECT 0.000000 1545.375000 2369.460000 1574.180000 ;
      RECT 1.100000 1544.475000 2369.460000 1545.375000 ;
      RECT 0.000000 1538.500000 2369.460000 1544.475000 ;
      RECT 0.000000 1537.600000 2368.360000 1538.500000 ;
      RECT 0.000000 1509.430000 2369.460000 1537.600000 ;
      RECT 1.100000 1508.530000 2369.460000 1509.430000 ;
      RECT 0.000000 1465.190000 2369.460000 1508.530000 ;
      RECT 0.000000 1464.290000 2368.360000 1465.190000 ;
      RECT 0.000000 1437.540000 2369.460000 1464.290000 ;
      RECT 1.100000 1436.640000 2369.460000 1437.540000 ;
      RECT 0.000000 1428.610000 2369.460000 1436.640000 ;
      RECT 0.000000 1427.710000 2368.360000 1428.610000 ;
      RECT 0.000000 1401.595000 2369.460000 1427.710000 ;
      RECT 1.100000 1400.695000 2369.460000 1401.595000 ;
      RECT 0.000000 1391.955000 2369.460000 1400.695000 ;
      RECT 0.000000 1391.055000 2368.360000 1391.955000 ;
      RECT 0.000000 1365.730000 2369.460000 1391.055000 ;
      RECT 1.100000 1364.830000 2369.460000 1365.730000 ;
      RECT 0.000000 1318.725000 2369.460000 1364.830000 ;
      RECT 0.000000 1317.825000 2368.360000 1318.725000 ;
      RECT 0.000000 1293.840000 2369.460000 1317.825000 ;
      RECT 1.100000 1292.940000 2369.460000 1293.840000 ;
      RECT 0.000000 1282.065000 2369.460000 1292.940000 ;
      RECT 0.000000 1281.165000 2368.360000 1282.065000 ;
      RECT 0.000000 1257.895000 2369.460000 1281.165000 ;
      RECT 1.100000 1256.995000 2369.460000 1257.895000 ;
      RECT 0.000000 1245.490000 2369.460000 1256.995000 ;
      RECT 0.000000 1244.590000 2368.360000 1245.490000 ;
      RECT 0.000000 1221.950000 2369.460000 1244.590000 ;
      RECT 1.100000 1221.050000 2369.460000 1221.950000 ;
      RECT 0.000000 1172.255000 2369.460000 1221.050000 ;
      RECT 0.000000 1171.355000 2368.360000 1172.255000 ;
      RECT 0.000000 1150.135000 2369.460000 1171.355000 ;
      RECT 1.100000 1149.235000 2369.460000 1150.135000 ;
      RECT 0.000000 1135.600000 2369.460000 1149.235000 ;
      RECT 0.000000 1134.700000 2368.360000 1135.600000 ;
      RECT 0.000000 1114.190000 2369.460000 1134.700000 ;
      RECT 1.100000 1113.290000 2369.460000 1114.190000 ;
      RECT 0.000000 1099.025000 2369.460000 1113.290000 ;
      RECT 0.000000 1098.125000 2368.360000 1099.025000 ;
      RECT 0.000000 1078.325000 2369.460000 1098.125000 ;
      RECT 1.100000 1077.425000 2369.460000 1078.325000 ;
      RECT 0.000000 1025.710000 2369.460000 1077.425000 ;
      RECT 0.000000 1024.810000 2368.360000 1025.710000 ;
      RECT 0.000000 1006.355000 2369.460000 1024.810000 ;
      RECT 1.100000 1005.455000 2369.460000 1006.355000 ;
      RECT 0.000000 989.135000 2369.460000 1005.455000 ;
      RECT 0.000000 988.235000 2368.360000 989.135000 ;
      RECT 0.000000 970.490000 2369.460000 988.235000 ;
      RECT 1.100000 969.590000 2369.460000 970.490000 ;
      RECT 0.000000 952.560000 2369.460000 969.590000 ;
      RECT 0.000000 951.660000 2368.360000 952.560000 ;
      RECT 0.000000 934.545000 2369.460000 951.660000 ;
      RECT 1.100000 933.645000 2369.460000 934.545000 ;
      RECT 0.000000 879.245000 2369.460000 933.645000 ;
      RECT 0.000000 878.345000 2368.360000 879.245000 ;
      RECT 0.000000 862.735000 2369.460000 878.345000 ;
      RECT 1.100000 861.835000 2369.460000 862.735000 ;
      RECT 0.000000 842.670000 2369.460000 861.835000 ;
      RECT 0.000000 841.770000 2368.360000 842.670000 ;
      RECT 0.000000 826.710000 2369.460000 841.770000 ;
      RECT 1.100000 825.810000 2369.460000 826.710000 ;
      RECT 0.000000 806.015000 2369.460000 825.810000 ;
      RECT 0.000000 805.115000 2368.360000 806.015000 ;
      RECT 0.000000 790.845000 2369.460000 805.115000 ;
      RECT 1.100000 789.945000 2369.460000 790.845000 ;
      RECT 0.000000 732.780000 2369.460000 789.945000 ;
      RECT 0.000000 731.880000 2368.360000 732.780000 ;
      RECT 0.000000 718.955000 2369.460000 731.880000 ;
      RECT 1.100000 718.055000 2369.460000 718.955000 ;
      RECT 0.000000 696.125000 2369.460000 718.055000 ;
      RECT 0.000000 695.225000 2368.360000 696.125000 ;
      RECT 0.000000 683.090000 2369.460000 695.225000 ;
      RECT 1.100000 682.190000 2369.460000 683.090000 ;
      RECT 0.000000 659.545000 2369.460000 682.190000 ;
      RECT 0.000000 658.645000 2368.360000 659.545000 ;
      RECT 0.000000 647.145000 2369.460000 658.645000 ;
      RECT 1.100000 646.245000 2369.460000 647.145000 ;
      RECT 0.000000 622.970000 2369.460000 646.245000 ;
      RECT 0.000000 622.070000 2368.360000 622.970000 ;
      RECT 0.000000 586.315000 2369.460000 622.070000 ;
      RECT 0.000000 585.415000 2368.360000 586.315000 ;
      RECT 0.000000 575.255000 2369.460000 585.415000 ;
      RECT 1.100000 574.355000 2369.460000 575.255000 ;
      RECT 0.000000 549.660000 2369.460000 574.355000 ;
      RECT 0.000000 548.760000 2368.360000 549.660000 ;
      RECT 0.000000 539.310000 2369.460000 548.760000 ;
      RECT 1.100000 538.410000 2369.460000 539.310000 ;
      RECT 0.000000 513.080000 2369.460000 538.410000 ;
      RECT 0.000000 512.180000 2368.360000 513.080000 ;
      RECT 0.000000 503.365000 2369.460000 512.180000 ;
      RECT 1.100000 502.465000 2369.460000 503.365000 ;
      RECT 0.000000 476.505000 2369.460000 502.465000 ;
      RECT 0.000000 475.605000 2368.360000 476.505000 ;
      RECT 0.000000 439.850000 2369.460000 475.605000 ;
      RECT 0.000000 438.950000 2368.360000 439.850000 ;
      RECT 0.000000 431.555000 2369.460000 438.950000 ;
      RECT 1.100000 430.655000 2369.460000 431.555000 ;
      RECT 0.000000 403.190000 2369.460000 430.655000 ;
      RECT 0.000000 402.290000 2368.360000 403.190000 ;
      RECT 0.000000 395.610000 2369.460000 402.290000 ;
      RECT 1.100000 394.710000 2369.460000 395.610000 ;
      RECT 0.000000 366.615000 2369.460000 394.710000 ;
      RECT 0.000000 365.715000 2368.360000 366.615000 ;
      RECT 0.000000 359.665000 2369.460000 365.715000 ;
      RECT 1.100000 358.765000 2369.460000 359.665000 ;
      RECT 0.000000 329.960000 2369.460000 358.765000 ;
      RECT 0.000000 329.060000 2368.360000 329.960000 ;
      RECT 0.000000 293.380000 2369.460000 329.060000 ;
      RECT 0.000000 292.480000 2368.360000 293.380000 ;
      RECT 0.000000 287.850000 2369.460000 292.480000 ;
      RECT 1.100000 286.950000 2369.460000 287.850000 ;
      RECT 0.000000 256.725000 2369.460000 286.950000 ;
      RECT 0.000000 255.825000 2368.360000 256.725000 ;
      RECT 0.000000 251.905000 2369.460000 255.825000 ;
      RECT 1.100000 251.005000 2369.460000 251.905000 ;
      RECT 0.000000 220.070000 2369.460000 251.005000 ;
      RECT 0.000000 219.170000 2368.360000 220.070000 ;
      RECT 0.000000 215.960000 2369.460000 219.170000 ;
      RECT 1.100000 215.060000 2369.460000 215.960000 ;
      RECT 0.000000 183.495000 2369.460000 215.060000 ;
      RECT 0.000000 182.595000 2368.360000 183.495000 ;
      RECT 0.000000 180.015000 2369.460000 182.595000 ;
      RECT 1.100000 179.115000 2369.460000 180.015000 ;
      RECT 0.000000 146.915000 2369.460000 179.115000 ;
      RECT 0.000000 146.015000 2368.360000 146.915000 ;
      RECT 0.000000 144.070000 2369.460000 146.015000 ;
      RECT 1.100000 143.170000 2369.460000 144.070000 ;
      RECT 0.000000 110.180000 2369.460000 143.170000 ;
      RECT 0.000000 109.280000 2368.360000 110.180000 ;
      RECT 0.000000 108.125000 2369.460000 109.280000 ;
      RECT 1.100000 107.225000 2369.460000 108.125000 ;
      RECT 0.000000 73.605000 2369.460000 107.225000 ;
      RECT 0.000000 72.705000 2368.360000 73.605000 ;
      RECT 0.000000 72.260000 2369.460000 72.705000 ;
      RECT 1.100000 71.360000 2369.460000 72.260000 ;
      RECT 0.000000 37.025000 2369.460000 71.360000 ;
      RECT 0.000000 36.125000 2368.360000 37.025000 ;
      RECT 0.000000 2.190000 2369.460000 36.125000 ;
      RECT 0.000000 1.290000 2368.360000 2.190000 ;
      RECT 0.000000 0.000000 2369.460000 1.290000 ;
    LAYER met4 ;
      RECT 0.000000 0.000000 2369.460000 2290.240000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
