magic
tech sky130A
magscale 1 2
timestamp 1647447581
<< metal1 >>
rect 56594 29860 56600 29912
rect 56652 29900 56658 29912
rect 57637 29900 57643 29912
rect 56652 29872 57643 29900
rect 56652 29860 56658 29872
rect 57637 29860 57643 29872
rect 57695 29860 57701 29912
rect 62114 29860 62120 29912
rect 62172 29900 62178 29912
rect 63094 29900 63100 29912
rect 62172 29872 63100 29900
rect 62172 29860 62178 29872
rect 63094 29860 63100 29872
rect 63152 29860 63158 29912
rect 71866 29792 71872 29844
rect 71924 29832 71930 29844
rect 73073 29832 73079 29844
rect 71924 29804 73079 29832
rect 71924 29792 71930 29804
rect 73073 29792 73079 29804
rect 73131 29792 73137 29844
rect 77294 29792 77300 29844
rect 77352 29832 77358 29844
rect 78547 29832 78553 29844
rect 77352 29804 78553 29832
rect 77352 29792 77358 29804
rect 78547 29792 78553 29804
rect 78605 29792 78611 29844
rect 80054 29792 80060 29844
rect 80112 29832 80118 29844
rect 81284 29832 81290 29844
rect 80112 29804 81290 29832
rect 80112 29792 80118 29804
rect 81284 29792 81290 29804
rect 81342 29792 81348 29844
rect 82814 29792 82820 29844
rect 82872 29832 82878 29844
rect 83987 29832 83993 29844
rect 82872 29804 83993 29832
rect 82872 29792 82878 29804
rect 83987 29792 83993 29804
rect 84045 29792 84051 29844
rect 85666 29792 85672 29844
rect 85724 29832 85730 29844
rect 86724 29832 86730 29844
rect 85724 29804 86730 29832
rect 85724 29792 85730 29804
rect 86724 29792 86730 29804
rect 86782 29792 86788 29844
rect 88426 29792 88432 29844
rect 88484 29832 88490 29844
rect 89444 29832 89450 29844
rect 88484 29804 89450 29832
rect 88484 29792 88490 29804
rect 89444 29792 89450 29804
rect 89502 29792 89508 29844
rect 111886 29792 111892 29844
rect 111944 29832 111950 29844
rect 113091 29832 113097 29844
rect 111944 29804 113097 29832
rect 111944 29792 111950 29804
rect 113091 29792 113097 29804
rect 113149 29792 113155 29844
rect 128354 29792 128360 29844
rect 128412 29832 128418 29844
rect 129479 29832 129485 29844
rect 128412 29804 129485 29832
rect 128412 29792 128418 29804
rect 129479 29792 129485 29804
rect 129537 29792 129543 29844
rect 133874 29792 133880 29844
rect 133932 29832 133938 29844
rect 134936 29832 134942 29844
rect 133932 29804 134942 29832
rect 133932 29792 133938 29804
rect 134936 29792 134942 29804
rect 134994 29792 135000 29844
rect 136634 29792 136640 29844
rect 136692 29832 136698 29844
rect 137673 29832 137679 29844
rect 136692 29804 137679 29832
rect 136692 29792 136698 29804
rect 137673 29792 137679 29804
rect 137731 29792 137737 29844
rect 139394 29792 139400 29844
rect 139452 29832 139458 29844
rect 140393 29832 140399 29844
rect 139452 29804 140399 29832
rect 139452 29792 139458 29804
rect 140393 29792 140399 29804
rect 140451 29792 140457 29844
rect 189074 29792 189080 29844
rect 189132 29832 189138 29844
rect 190407 29832 190413 29844
rect 189132 29804 190413 29832
rect 189132 29792 189138 29804
rect 190407 29792 190413 29804
rect 190465 29792 190471 29844
rect 197446 29792 197452 29844
rect 197504 29832 197510 29844
rect 198567 29832 198573 29844
rect 197504 29804 198573 29832
rect 197504 29792 197510 29804
rect 198567 29792 198573 29804
rect 198625 29792 198631 29844
rect 200114 29792 200120 29844
rect 200172 29832 200178 29844
rect 201304 29832 201310 29844
rect 200172 29804 201310 29832
rect 200172 29792 200178 29804
rect 201304 29792 201310 29804
rect 201362 29792 201368 29844
rect 205634 29792 205640 29844
rect 205692 29832 205698 29844
rect 206744 29832 206750 29844
rect 205692 29804 206750 29832
rect 205692 29792 205698 29804
rect 206744 29792 206750 29804
rect 206802 29792 206808 29844
rect 211154 29792 211160 29844
rect 211212 29832 211218 29844
rect 212235 29832 212241 29844
rect 211212 29804 212241 29832
rect 211212 29792 211218 29804
rect 212235 29792 212241 29804
rect 212293 29792 212299 29844
rect 231854 29792 231860 29844
rect 231912 29832 231918 29844
rect 233128 29832 233134 29844
rect 231912 29804 233134 29832
rect 231912 29792 231918 29804
rect 233128 29792 233134 29804
rect 233186 29792 233192 29844
rect 237374 29792 237380 29844
rect 237432 29832 237438 29844
rect 238602 29832 238608 29844
rect 237432 29804 238608 29832
rect 237432 29792 237438 29804
rect 238602 29792 238608 29804
rect 238660 29792 238666 29844
rect 240134 29792 240140 29844
rect 240192 29832 240198 29844
rect 241356 29832 241362 29844
rect 240192 29804 241362 29832
rect 240192 29792 240198 29804
rect 241356 29792 241362 29804
rect 241414 29792 241420 29844
rect 242894 29792 242900 29844
rect 242952 29832 242958 29844
rect 244042 29832 244048 29844
rect 242952 29804 244048 29832
rect 242952 29792 242958 29804
rect 244042 29792 244048 29804
rect 244100 29792 244106 29844
rect 259454 29792 259460 29844
rect 259512 29832 259518 29844
rect 260430 29832 260436 29844
rect 259512 29804 260436 29832
rect 259512 29792 259518 29804
rect 260430 29792 260436 29804
rect 260488 29792 260494 29844
rect 274634 29792 274640 29844
rect 274692 29832 274698 29844
rect 275883 29832 275889 29844
rect 274692 29804 275889 29832
rect 274692 29792 274698 29804
rect 275883 29792 275889 29804
rect 275941 29792 275947 29844
rect 277486 29792 277492 29844
rect 277544 29832 277550 29844
rect 278603 29832 278609 29844
rect 277544 29804 278609 29832
rect 277544 29792 277550 29804
rect 278603 29792 278609 29804
rect 278661 29792 278667 29844
rect 285674 29792 285680 29844
rect 285732 29832 285738 29844
rect 286831 29832 286837 29844
rect 285732 29804 286837 29832
rect 285732 29792 285738 29804
rect 286831 29792 286837 29804
rect 286889 29792 286895 29844
rect 291194 29792 291200 29844
rect 291252 29832 291258 29844
rect 292254 29832 292260 29844
rect 291252 29804 292260 29832
rect 291252 29792 291258 29804
rect 292254 29792 292260 29804
rect 292312 29792 292318 29844
rect 311894 29792 311900 29844
rect 311952 29832 311958 29844
rect 313147 29832 313153 29844
rect 311952 29804 313153 29832
rect 311952 29792 311958 29804
rect 313147 29792 313153 29804
rect 313205 29792 313211 29844
rect 314746 29792 314752 29844
rect 314804 29832 314810 29844
rect 315884 29832 315890 29844
rect 314804 29804 315890 29832
rect 314804 29792 314810 29804
rect 315884 29792 315890 29804
rect 315942 29792 315948 29844
rect 317414 29792 317420 29844
rect 317472 29832 317478 29844
rect 318621 29832 318627 29844
rect 317472 29804 318627 29832
rect 317472 29792 317478 29804
rect 318621 29792 318627 29804
rect 318679 29792 318685 29844
rect 346394 29792 346400 29844
rect 346452 29832 346458 29844
rect 347725 29832 347731 29844
rect 346452 29804 347731 29832
rect 346452 29792 346458 29804
rect 347725 29792 347731 29804
rect 347783 29792 347789 29844
rect 352006 29792 352012 29844
rect 352064 29832 352070 29844
rect 353182 29832 353188 29844
rect 352064 29804 353188 29832
rect 352064 29792 352070 29804
rect 353182 29792 353188 29804
rect 353240 29792 353246 29844
rect 357434 29792 357440 29844
rect 357492 29832 357498 29844
rect 358639 29832 358645 29844
rect 357492 29804 358645 29832
rect 357492 29792 357498 29804
rect 358639 29792 358645 29804
rect 358697 29792 358703 29844
rect 362954 29792 362960 29844
rect 363012 29832 363018 29844
rect 364096 29832 364102 29844
rect 363012 29804 364102 29832
rect 363012 29792 363018 29804
rect 364096 29792 364102 29804
rect 364154 29792 364160 29844
rect 373994 29792 374000 29844
rect 374052 29832 374058 29844
rect 375010 29832 375016 29844
rect 374052 29804 375016 29832
rect 374052 29792 374058 29804
rect 375010 29792 375016 29804
rect 375068 29792 375074 29844
rect 389174 29792 389180 29844
rect 389232 29832 389238 29844
rect 390463 29832 390469 29844
rect 389232 29804 390469 29832
rect 389232 29792 389238 29804
rect 390463 29792 390469 29804
rect 390521 29792 390527 29844
rect 405734 29792 405740 29844
rect 405792 29832 405798 29844
rect 406851 29832 406857 29844
rect 405792 29804 406857 29832
rect 405792 29792 405798 29804
rect 406851 29792 406857 29804
rect 406909 29792 406915 29844
rect 426526 29792 426532 29844
rect 426584 29832 426590 29844
rect 427744 29832 427750 29844
rect 426584 29804 427750 29832
rect 426584 29792 426590 29804
rect 427744 29792 427750 29804
rect 427802 29792 427808 29844
rect 431954 29792 431960 29844
rect 432012 29832 432018 29844
rect 433167 29832 433173 29844
rect 432012 29804 433173 29832
rect 432012 29792 432018 29804
rect 433167 29792 433173 29804
rect 433225 29792 433231 29844
rect 434806 29792 434812 29844
rect 434864 29832 434870 29844
rect 435921 29832 435927 29844
rect 434864 29804 435927 29832
rect 434864 29792 434870 29804
rect 435921 29792 435927 29804
rect 435979 29792 435985 29844
rect 448514 29792 448520 29844
rect 448572 29832 448578 29844
rect 449572 29832 449578 29844
rect 448572 29804 449578 29832
rect 448572 29792 448578 29804
rect 449572 29792 449578 29804
rect 449630 29792 449636 29844
rect 474826 29792 474832 29844
rect 474884 29832 474890 29844
rect 475973 29832 475979 29844
rect 474884 29804 475979 29832
rect 474884 29792 474890 29804
rect 475973 29792 475979 29804
rect 476031 29792 476037 29844
rect 488534 29792 488540 29844
rect 488592 29832 488598 29844
rect 489607 29832 489613 29844
rect 488592 29804 489613 29832
rect 488592 29792 488598 29804
rect 489607 29792 489613 29804
rect 489665 29792 489671 29844
rect 491294 29792 491300 29844
rect 491352 29832 491358 29844
rect 492310 29832 492316 29844
rect 491352 29804 492316 29832
rect 491352 29792 491358 29804
rect 492310 29792 492316 29804
rect 492368 29792 492374 29844
rect 494054 29792 494060 29844
rect 494112 29832 494118 29844
rect 495047 29832 495053 29844
rect 494112 29804 495053 29832
rect 494112 29792 494118 29804
rect 495047 29792 495053 29804
rect 495105 29792 495111 29844
rect 201494 28500 201500 28552
rect 201552 28540 201558 28552
rect 403158 28540 403164 28552
rect 201552 28512 403164 28540
rect 201552 28500 201558 28512
rect 403158 28500 403164 28512
rect 403216 28500 403222 28552
rect 194594 28432 194600 28484
rect 194652 28472 194658 28484
rect 401410 28472 401416 28484
rect 194652 28444 401416 28472
rect 194652 28432 194658 28444
rect 401410 28432 401416 28444
rect 401468 28432 401474 28484
rect 185026 28364 185032 28416
rect 185084 28404 185090 28416
rect 398650 28404 398656 28416
rect 185084 28376 398656 28404
rect 185084 28364 185090 28376
rect 398650 28364 398656 28376
rect 398708 28364 398714 28416
rect 176654 28296 176660 28348
rect 176712 28336 176718 28348
rect 396810 28336 396816 28348
rect 176712 28308 396816 28336
rect 176712 28296 176718 28308
rect 396810 28296 396816 28308
rect 396868 28296 396874 28348
rect 162854 28228 162860 28280
rect 162912 28268 162918 28280
rect 393222 28268 393228 28280
rect 162912 28240 393228 28268
rect 162912 28228 162918 28240
rect 393222 28228 393228 28240
rect 393280 28228 393286 28280
rect 64874 28092 64880 28144
rect 64932 28132 64938 28144
rect 65794 28132 65800 28144
rect 64932 28104 65800 28132
rect 64932 28092 64938 28104
rect 65794 28092 65800 28104
rect 65852 28092 65858 28144
rect 67634 28092 67640 28144
rect 67692 28132 67698 28144
rect 68554 28132 68560 28144
rect 67692 28104 68560 28132
rect 67692 28092 67698 28104
rect 68554 28092 68560 28104
rect 68612 28092 68618 28144
rect 102134 28092 102140 28144
rect 102192 28132 102198 28144
rect 103054 28132 103060 28144
rect 102192 28104 103060 28132
rect 102192 28092 102198 28104
rect 103054 28092 103060 28104
rect 103112 28092 103118 28144
rect 104894 28092 104900 28144
rect 104952 28132 104958 28144
rect 105814 28132 105820 28144
rect 104952 28104 105820 28132
rect 104952 28092 104958 28104
rect 105814 28092 105820 28104
rect 105872 28092 105878 28144
rect 110414 28092 110420 28144
rect 110472 28132 110478 28144
rect 111242 28132 111248 28144
rect 110472 28104 111248 28132
rect 110472 28092 110478 28104
rect 111242 28092 111248 28104
rect 111300 28092 111306 28144
rect 114646 28092 114652 28144
rect 114704 28132 114710 28144
rect 115842 28132 115848 28144
rect 114704 28104 115848 28132
rect 114704 28092 114710 28104
rect 115842 28092 115848 28104
rect 115900 28092 115906 28144
rect 142154 28092 142160 28144
rect 142212 28132 142218 28144
rect 143074 28132 143080 28144
rect 142212 28104 143080 28132
rect 142212 28092 142218 28104
rect 143074 28092 143080 28104
rect 143132 28092 143138 28144
rect 147674 28092 147680 28144
rect 147732 28132 147738 28144
rect 148502 28132 148508 28144
rect 147732 28104 148508 28132
rect 147732 28092 147738 28104
rect 148502 28092 148508 28104
rect 148560 28092 148566 28144
rect 151906 28092 151912 28144
rect 151964 28132 151970 28144
rect 153102 28132 153108 28144
rect 151964 28104 153108 28132
rect 151964 28092 151970 28104
rect 153102 28092 153108 28104
rect 153160 28092 153166 28144
rect 182174 28092 182180 28144
rect 182232 28132 182238 28144
rect 183094 28132 183100 28144
rect 182232 28104 183100 28132
rect 182232 28092 182238 28104
rect 183094 28092 183100 28104
rect 183152 28092 183158 28144
rect 222194 28092 222200 28144
rect 222252 28132 222258 28144
rect 223114 28132 223120 28144
rect 222252 28104 223120 28132
rect 222252 28092 222258 28104
rect 223114 28092 223120 28104
rect 223172 28092 223178 28144
rect 269206 28092 269212 28144
rect 269264 28132 269270 28144
rect 270402 28132 270408 28144
rect 269264 28104 270408 28132
rect 269264 28092 269270 28104
rect 270402 28092 270408 28104
rect 270460 28092 270466 28144
rect 302234 28092 302240 28144
rect 302292 28132 302298 28144
rect 303154 28132 303160 28144
rect 302292 28104 303160 28132
rect 302292 28092 302298 28104
rect 303154 28092 303160 28104
rect 303212 28092 303218 28144
rect 309226 28092 309232 28144
rect 309284 28132 309290 28144
rect 310422 28132 310428 28144
rect 309284 28104 310428 28132
rect 309284 28092 309290 28104
rect 310422 28092 310428 28104
rect 310480 28092 310486 28144
rect 339494 28092 339500 28144
rect 339552 28132 339558 28144
rect 340414 28132 340420 28144
rect 339552 28104 340420 28132
rect 339552 28092 339558 28104
rect 340414 28092 340420 28104
rect 340472 28092 340478 28144
rect 429286 28092 429292 28144
rect 429344 28132 429350 28144
rect 430482 28132 430488 28144
rect 429344 28104 430488 28132
rect 429344 28092 429350 28104
rect 430482 28092 430488 28104
rect 430540 28092 430546 28144
rect 456794 28092 456800 28144
rect 456852 28132 456858 28144
rect 457714 28132 457720 28144
rect 456852 28104 457720 28132
rect 456852 28092 456858 28104
rect 457714 28092 457720 28104
rect 457772 28092 457778 28144
rect 459554 28092 459560 28144
rect 459612 28132 459618 28144
rect 460474 28132 460480 28144
rect 459612 28104 460480 28132
rect 459612 28092 459618 28104
rect 460474 28092 460480 28104
rect 460532 28092 460538 28144
rect 69014 27548 69020 27600
rect 69072 27588 69078 27600
rect 72142 27588 72148 27600
rect 69072 27560 72148 27588
rect 69072 27548 69078 27560
rect 72142 27548 72148 27560
rect 72200 27548 72206 27600
rect 90358 27548 90364 27600
rect 90416 27588 90422 27600
rect 92198 27588 92204 27600
rect 90416 27560 92204 27588
rect 90416 27548 90422 27560
rect 92198 27548 92204 27560
rect 92256 27548 92262 27600
rect 106918 27548 106924 27600
rect 106976 27588 106982 27600
rect 107654 27588 107660 27600
rect 106976 27560 107660 27588
rect 106976 27548 106982 27560
rect 107654 27548 107660 27560
rect 107712 27548 107718 27600
rect 108942 27548 108948 27600
rect 109000 27588 109006 27600
rect 109494 27588 109500 27600
rect 109000 27560 109500 27588
rect 109000 27548 109006 27560
rect 109494 27548 109500 27560
rect 109552 27548 109558 27600
rect 114002 27548 114008 27600
rect 114060 27588 114066 27600
rect 115934 27588 115940 27600
rect 114060 27560 115940 27588
rect 114060 27548 114066 27560
rect 115934 27548 115940 27560
rect 115992 27548 115998 27600
rect 117222 27548 117228 27600
rect 117280 27588 117286 27600
rect 117682 27588 117688 27600
rect 117280 27560 117688 27588
rect 117280 27548 117286 27560
rect 117682 27548 117688 27560
rect 117740 27548 117746 27600
rect 126238 27548 126244 27600
rect 126296 27588 126302 27600
rect 127618 27588 127624 27600
rect 126296 27560 127624 27588
rect 126296 27548 126302 27560
rect 127618 27548 127624 27560
rect 127676 27548 127682 27600
rect 155218 27548 155224 27600
rect 155276 27588 155282 27600
rect 158530 27588 158536 27600
rect 155276 27560 158536 27588
rect 155276 27548 155282 27560
rect 158530 27548 158536 27560
rect 158588 27548 158594 27600
rect 163130 27548 163136 27600
rect 163188 27588 163194 27600
rect 170398 27588 170404 27600
rect 163188 27560 170404 27588
rect 163188 27548 163194 27560
rect 170398 27548 170404 27560
rect 170456 27548 170462 27600
rect 171318 27548 171324 27600
rect 171376 27588 171382 27600
rect 173158 27588 173164 27600
rect 171376 27560 173164 27588
rect 171376 27548 171382 27560
rect 173158 27548 173164 27560
rect 173216 27548 173222 27600
rect 185854 27548 185860 27600
rect 185912 27588 185918 27600
rect 186958 27588 186964 27600
rect 185912 27560 186964 27588
rect 185912 27548 185918 27560
rect 186958 27548 186964 27560
rect 187016 27548 187022 27600
rect 204070 27548 204076 27600
rect 204128 27588 204134 27600
rect 205542 27588 205548 27600
rect 204128 27560 205548 27588
rect 204128 27548 204134 27560
rect 205542 27548 205548 27560
rect 205600 27548 205606 27600
rect 243170 27548 243176 27600
rect 243228 27588 243234 27600
rect 244918 27588 244924 27600
rect 243228 27560 244924 27588
rect 243228 27548 243234 27560
rect 244918 27548 244924 27560
rect 244976 27548 244982 27600
rect 254026 27548 254032 27600
rect 254084 27588 254090 27600
rect 256602 27588 256608 27600
rect 254084 27560 256608 27588
rect 254084 27548 254090 27560
rect 256602 27548 256608 27560
rect 256660 27548 256666 27600
rect 264974 27548 264980 27600
rect 265032 27588 265038 27600
rect 267642 27588 267648 27600
rect 265032 27560 267648 27588
rect 265032 27548 265038 27560
rect 267642 27548 267648 27560
rect 267700 27548 267706 27600
rect 282178 27548 282184 27600
rect 282236 27588 282242 27600
rect 283190 27588 283196 27600
rect 282236 27560 283196 27588
rect 282236 27548 282242 27560
rect 283190 27548 283196 27560
rect 283248 27548 283254 27600
rect 300118 27548 300124 27600
rect 300176 27588 300182 27600
rect 301314 27588 301320 27600
rect 300176 27560 301320 27588
rect 300176 27548 300182 27560
rect 301314 27548 301320 27560
rect 301372 27548 301378 27600
rect 313918 27548 313924 27600
rect 313976 27588 313982 27600
rect 314930 27588 314936 27600
rect 313976 27560 314936 27588
rect 313976 27548 313982 27560
rect 314930 27548 314936 27560
rect 314988 27548 314994 27600
rect 325878 27548 325884 27600
rect 325936 27588 325942 27600
rect 327718 27588 327724 27600
rect 325936 27560 327724 27588
rect 325936 27548 325942 27560
rect 327718 27548 327724 27560
rect 327776 27548 327782 27600
rect 355962 27548 355968 27600
rect 356020 27588 356026 27600
rect 356698 27588 356704 27600
rect 356020 27560 356704 27588
rect 356020 27548 356026 27560
rect 356698 27548 356704 27560
rect 356756 27548 356762 27600
rect 396718 27548 396724 27600
rect 396776 27588 396782 27600
rect 397730 27588 397736 27600
rect 396776 27560 397736 27588
rect 396776 27548 396782 27560
rect 397730 27548 397736 27560
rect 397788 27548 397794 27600
rect 407758 27548 407764 27600
rect 407816 27588 407822 27600
rect 408678 27588 408684 27600
rect 407816 27560 408684 27588
rect 407816 27548 407822 27560
rect 408678 27548 408684 27560
rect 408736 27548 408742 27600
rect 416682 27548 416688 27600
rect 416740 27588 416746 27600
rect 421282 27588 421288 27600
rect 416740 27560 421288 27588
rect 416740 27548 416746 27560
rect 421282 27548 421288 27560
rect 421340 27548 421346 27600
rect 425698 27548 425704 27600
rect 425756 27588 425762 27600
rect 428642 27588 428648 27600
rect 425756 27560 428648 27588
rect 425756 27548 425762 27560
rect 428642 27548 428648 27560
rect 428700 27548 428706 27600
rect 465258 27548 465264 27600
rect 465316 27588 465322 27600
rect 470502 27588 470508 27600
rect 465316 27560 470508 27588
rect 465316 27548 465322 27560
rect 470502 27548 470508 27560
rect 470560 27548 470566 27600
rect 473262 27548 473268 27600
rect 473320 27588 473326 27600
rect 474734 27588 474740 27600
rect 473320 27560 474740 27588
rect 473320 27548 473326 27560
rect 474734 27548 474740 27560
rect 474792 27548 474798 27600
rect 481358 27548 481364 27600
rect 481416 27588 481422 27600
rect 485038 27588 485044 27600
rect 481416 27560 485044 27588
rect 481416 27548 481422 27560
rect 485038 27548 485044 27560
rect 485096 27548 485102 27600
rect 109034 27480 109040 27532
rect 109092 27520 109098 27532
rect 112162 27520 112168 27532
rect 109092 27492 112168 27520
rect 109092 27480 109098 27492
rect 112162 27480 112168 27492
rect 112220 27480 112226 27532
rect 225874 27480 225880 27532
rect 225932 27520 225938 27532
rect 249058 27520 249064 27532
rect 225932 27492 249064 27520
rect 225932 27480 225938 27492
rect 249058 27480 249064 27492
rect 249116 27480 249122 27532
rect 298738 27480 298744 27532
rect 298796 27520 298802 27532
rect 300394 27520 300400 27532
rect 298796 27492 300400 27520
rect 298796 27480 298802 27492
rect 300394 27480 300400 27492
rect 300452 27480 300458 27532
rect 361390 27480 361396 27532
rect 361448 27520 361454 27532
rect 376110 27520 376116 27532
rect 361448 27492 376116 27520
rect 361448 27480 361454 27492
rect 376110 27480 376116 27492
rect 376168 27480 376174 27532
rect 461026 27480 461032 27532
rect 461084 27520 461090 27532
rect 469582 27520 469588 27532
rect 461084 27492 469588 27520
rect 461084 27480 461090 27492
rect 469582 27480 469588 27492
rect 469640 27480 469646 27532
rect 214926 27412 214932 27464
rect 214984 27452 214990 27464
rect 273898 27452 273904 27464
rect 214984 27424 273904 27452
rect 214984 27412 214990 27424
rect 273898 27412 273904 27424
rect 273956 27412 273962 27464
rect 368658 27412 368664 27464
rect 368716 27452 368722 27464
rect 414658 27452 414664 27464
rect 368716 27424 414664 27452
rect 368716 27412 368722 27424
rect 414658 27412 414664 27424
rect 414716 27412 414722 27464
rect 207658 27344 207664 27396
rect 207716 27384 207722 27396
rect 291838 27384 291844 27396
rect 207716 27356 291844 27384
rect 207716 27344 207722 27356
rect 291838 27344 291844 27356
rect 291896 27344 291902 27396
rect 336826 27344 336832 27396
rect 336884 27384 336890 27396
rect 353386 27384 353392 27396
rect 336884 27356 353392 27384
rect 336884 27344 336890 27356
rect 353386 27344 353392 27356
rect 353444 27344 353450 27396
rect 362310 27344 362316 27396
rect 362368 27384 362374 27396
rect 410518 27384 410524 27396
rect 362368 27356 410524 27384
rect 362368 27344 362374 27356
rect 410518 27344 410524 27356
rect 410576 27344 410582 27396
rect 413278 27344 413284 27396
rect 413336 27384 413342 27396
rect 426802 27384 426808 27396
rect 413336 27356 426808 27384
rect 413336 27344 413342 27356
rect 426802 27344 426808 27356
rect 426860 27344 426866 27396
rect 203150 27276 203156 27328
rect 203208 27316 203214 27328
rect 296070 27316 296076 27328
rect 203208 27288 296076 27316
rect 203208 27276 203214 27288
rect 296070 27276 296076 27288
rect 296128 27276 296134 27328
rect 348602 27276 348608 27328
rect 348660 27316 348666 27328
rect 364978 27316 364984 27328
rect 348660 27288 364984 27316
rect 348660 27276 348666 27288
rect 364978 27276 364984 27288
rect 365036 27276 365042 27328
rect 367738 27276 367744 27328
rect 367796 27316 367802 27328
rect 419534 27316 419540 27328
rect 367796 27288 419540 27316
rect 367796 27276 367802 27288
rect 419534 27276 419540 27288
rect 419592 27276 419598 27328
rect 454034 27276 454040 27328
rect 454092 27316 454098 27328
rect 467742 27316 467748 27328
rect 454092 27288 467748 27316
rect 454092 27276 454098 27288
rect 467742 27276 467748 27288
rect 467800 27276 467806 27328
rect 95142 27208 95148 27260
rect 95200 27248 95206 27260
rect 95786 27248 95792 27260
rect 95200 27220 95792 27248
rect 95200 27208 95206 27220
rect 95786 27208 95792 27220
rect 95844 27208 95850 27260
rect 219526 27208 219532 27260
rect 219584 27248 219590 27260
rect 339126 27248 339132 27260
rect 219584 27220 339132 27248
rect 219584 27208 219590 27220
rect 339126 27208 339132 27220
rect 339184 27208 339190 27260
rect 341334 27208 341340 27260
rect 341392 27248 341398 27260
rect 360470 27248 360476 27260
rect 341392 27220 360476 27248
rect 341392 27208 341398 27220
rect 360470 27208 360476 27220
rect 360528 27208 360534 27260
rect 380434 27208 380440 27260
rect 380492 27248 380498 27260
rect 453298 27248 453304 27260
rect 380492 27220 453304 27248
rect 380492 27208 380498 27220
rect 453298 27208 453304 27220
rect 453356 27208 453362 27260
rect 130378 27140 130384 27192
rect 130436 27180 130442 27192
rect 131298 27180 131304 27192
rect 130436 27152 131304 27180
rect 130436 27140 130442 27152
rect 131298 27140 131304 27152
rect 131356 27140 131362 27192
rect 196802 27140 196808 27192
rect 196860 27180 196866 27192
rect 242158 27180 242164 27192
rect 196860 27152 242164 27180
rect 196860 27140 196866 27152
rect 242158 27140 242164 27152
rect 242216 27140 242222 27192
rect 261386 27140 261392 27192
rect 261444 27180 261450 27192
rect 407850 27180 407856 27192
rect 261444 27152 407856 27180
rect 261444 27140 261450 27152
rect 407850 27140 407856 27152
rect 407908 27140 407914 27192
rect 410426 27140 410432 27192
rect 410484 27180 410490 27192
rect 415946 27180 415952 27192
rect 410484 27152 415952 27180
rect 410484 27140 410490 27152
rect 415946 27140 415952 27152
rect 416004 27140 416010 27192
rect 418798 27140 418804 27192
rect 418856 27180 418862 27192
rect 440418 27180 440424 27192
rect 418856 27152 440424 27180
rect 418856 27140 418862 27152
rect 440418 27140 440424 27152
rect 440476 27140 440482 27192
rect 449894 27140 449900 27192
rect 449952 27180 449958 27192
rect 466822 27180 466828 27192
rect 449952 27152 466828 27180
rect 449952 27140 449958 27152
rect 466822 27140 466828 27152
rect 466880 27140 466886 27192
rect 184934 27072 184940 27124
rect 184992 27112 184998 27124
rect 246298 27112 246304 27124
rect 184992 27084 246304 27112
rect 184992 27072 184998 27084
rect 246298 27072 246304 27084
rect 246356 27072 246362 27124
rect 249518 27072 249524 27124
rect 249576 27112 249582 27124
rect 396810 27112 396816 27124
rect 249576 27084 396816 27112
rect 249576 27072 249582 27084
rect 396810 27072 396816 27084
rect 396868 27072 396874 27124
rect 403618 27072 403624 27124
rect 403676 27112 403682 27124
rect 437750 27112 437756 27124
rect 403676 27084 437756 27112
rect 403676 27072 403682 27084
rect 437750 27072 437756 27084
rect 437808 27072 437814 27124
rect 447226 27072 447232 27124
rect 447284 27112 447290 27124
rect 465994 27112 466000 27124
rect 447284 27084 466000 27112
rect 447284 27072 447290 27084
rect 465994 27072 466000 27084
rect 466052 27072 466058 27124
rect 480438 27072 480444 27124
rect 480496 27112 480502 27124
rect 503714 27112 503720 27124
rect 480496 27084 503720 27112
rect 480496 27072 480502 27084
rect 503714 27072 503720 27084
rect 503772 27072 503778 27124
rect 143534 27004 143540 27056
rect 143592 27044 143598 27056
rect 155862 27044 155868 27056
rect 143592 27016 155868 27044
rect 143592 27004 143598 27016
rect 155862 27004 155868 27016
rect 155920 27004 155926 27056
rect 166810 27004 166816 27056
rect 166868 27044 166874 27056
rect 184198 27044 184204 27056
rect 166868 27016 184204 27044
rect 166868 27004 166874 27016
rect 184198 27004 184204 27016
rect 184256 27004 184262 27056
rect 189442 27004 189448 27056
rect 189500 27044 189506 27056
rect 199378 27044 199384 27056
rect 189500 27016 199384 27044
rect 189500 27004 189506 27016
rect 199378 27004 199384 27016
rect 199436 27004 199442 27056
rect 240410 27004 240416 27056
rect 240468 27044 240474 27056
rect 418890 27044 418896 27056
rect 240468 27016 418896 27044
rect 240468 27004 240474 27016
rect 418890 27004 418896 27016
rect 418948 27004 418954 27056
rect 421558 27004 421564 27056
rect 421616 27044 421622 27056
rect 425882 27044 425888 27056
rect 421616 27016 425888 27044
rect 421616 27004 421622 27016
rect 425882 27004 425888 27016
rect 425940 27004 425946 27056
rect 440234 27004 440240 27056
rect 440292 27044 440298 27056
rect 464154 27044 464160 27056
rect 440292 27016 464160 27044
rect 440292 27004 440298 27016
rect 464154 27004 464160 27016
rect 464212 27004 464218 27056
rect 485958 27004 485964 27056
rect 486016 27044 486022 27056
rect 512638 27044 512644 27056
rect 486016 27016 512644 27044
rect 486016 27004 486022 27016
rect 512638 27004 512644 27016
rect 512696 27004 512702 27056
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 145834 26976 145840 26988
rect 15896 26948 145840 26976
rect 15896 26936 15902 26948
rect 145834 26936 145840 26948
rect 145892 26936 145898 26988
rect 146294 26936 146300 26988
rect 146352 26976 146358 26988
rect 156782 26976 156788 26988
rect 146352 26948 156788 26976
rect 146352 26936 146358 26948
rect 156782 26936 156788 26948
rect 156840 26936 156846 26988
rect 172238 26936 172244 26988
rect 172296 26976 172302 26988
rect 191098 26976 191104 26988
rect 172296 26948 191104 26976
rect 172296 26936 172302 26948
rect 191098 26936 191104 26948
rect 191156 26936 191162 26988
rect 191926 26936 191932 26988
rect 191984 26976 191990 26988
rect 193122 26976 193128 26988
rect 191984 26948 193128 26976
rect 191984 26936 191990 26948
rect 193122 26936 193128 26948
rect 193180 26936 193186 26988
rect 242250 26936 242256 26988
rect 242308 26976 242314 26988
rect 424318 26976 424324 26988
rect 242308 26948 424324 26976
rect 242308 26936 242314 26948
rect 424318 26936 424324 26948
rect 424376 26936 424382 26988
rect 424410 26936 424416 26988
rect 424468 26976 424474 26988
rect 434990 26976 434996 26988
rect 424468 26948 434996 26976
rect 424468 26936 424474 26948
rect 434990 26936 434996 26948
rect 435048 26936 435054 26988
rect 436094 26936 436100 26988
rect 436152 26976 436158 26988
rect 463234 26976 463240 26988
rect 436152 26948 463240 26976
rect 436152 26936 436158 26948
rect 463234 26936 463240 26948
rect 463292 26936 463298 26988
rect 482278 26936 482284 26988
rect 482336 26976 482342 26988
rect 510614 26976 510620 26988
rect 482336 26948 510620 26976
rect 482336 26936 482342 26948
rect 510614 26936 510620 26948
rect 510672 26936 510678 26988
rect 10318 26868 10324 26920
rect 10376 26908 10382 26920
rect 149514 26908 149520 26920
rect 10376 26880 149520 26908
rect 10376 26868 10382 26880
rect 149514 26868 149520 26880
rect 149572 26868 149578 26920
rect 150434 26868 150440 26920
rect 150492 26908 150498 26920
rect 157702 26908 157708 26920
rect 150492 26880 157708 26908
rect 150492 26868 150498 26880
rect 157702 26868 157708 26880
rect 157760 26868 157766 26920
rect 161290 26868 161296 26920
rect 161348 26908 161354 26920
rect 164234 26908 164240 26920
rect 161348 26880 164240 26908
rect 161348 26868 161354 26880
rect 164234 26868 164240 26880
rect 164292 26868 164298 26920
rect 167638 26868 167644 26920
rect 167696 26908 167702 26920
rect 175918 26908 175924 26920
rect 167696 26880 175924 26908
rect 167696 26868 167702 26880
rect 175918 26868 175924 26880
rect 175976 26868 175982 26920
rect 176746 26868 176752 26920
rect 176804 26908 176810 26920
rect 224218 26908 224224 26920
rect 176804 26880 224224 26908
rect 176804 26868 176810 26880
rect 224218 26868 224224 26880
rect 224276 26868 224282 26920
rect 230382 26868 230388 26920
rect 230440 26908 230446 26920
rect 428458 26908 428464 26920
rect 230440 26880 428464 26908
rect 230440 26868 230446 26880
rect 428458 26868 428464 26880
rect 428516 26868 428522 26920
rect 429378 26868 429384 26920
rect 429436 26908 429442 26920
rect 461394 26908 461400 26920
rect 429436 26880 461400 26908
rect 429436 26868 429442 26880
rect 461394 26868 461400 26880
rect 461452 26868 461458 26920
rect 477770 26868 477776 26920
rect 477828 26908 477834 26920
rect 492674 26908 492680 26920
rect 477828 26880 492680 26908
rect 477828 26868 477834 26880
rect 492674 26868 492680 26880
rect 492732 26868 492738 26920
rect 500494 26868 500500 26920
rect 500552 26908 500558 26920
rect 569218 26908 569224 26920
rect 500552 26880 569224 26908
rect 500552 26868 500558 26880
rect 569218 26868 569224 26880
rect 569276 26868 569282 26920
rect 271966 26800 271972 26852
rect 272024 26840 272030 26852
rect 273162 26840 273168 26852
rect 272024 26812 273168 26840
rect 272024 26800 272030 26812
rect 273162 26800 273168 26812
rect 273220 26800 273226 26852
rect 157518 26664 157524 26716
rect 157576 26704 157582 26716
rect 159450 26704 159456 26716
rect 157576 26676 159456 26704
rect 157576 26664 157582 26676
rect 159450 26664 159456 26676
rect 159508 26664 159514 26716
rect 77662 26324 77668 26376
rect 77720 26364 77726 26376
rect 79318 26364 79324 26376
rect 77720 26336 79324 26364
rect 77720 26324 77726 26336
rect 79318 26324 79324 26336
rect 79376 26324 79382 26376
rect 93118 26324 93124 26376
rect 93176 26364 93182 26376
rect 94038 26364 94044 26376
rect 93176 26336 94044 26364
rect 93176 26324 93182 26336
rect 94038 26324 94044 26336
rect 94096 26324 94102 26376
rect 296806 26364 296812 26376
rect 296686 26336 296812 26364
rect 54478 26256 54484 26308
rect 54536 26296 54542 26308
rect 55858 26296 55864 26308
rect 54536 26268 55864 26296
rect 54536 26256 54542 26268
rect 55858 26256 55864 26268
rect 55916 26256 55922 26308
rect 74074 26256 74080 26308
rect 74132 26296 74138 26308
rect 75914 26296 75920 26308
rect 74132 26268 75920 26296
rect 74132 26256 74138 26268
rect 75914 26256 75920 26268
rect 75972 26256 75978 26308
rect 295978 26256 295984 26308
rect 296036 26296 296042 26308
rect 296686 26296 296714 26336
rect 296806 26324 296812 26336
rect 296864 26324 296870 26376
rect 379606 26324 379612 26376
rect 379664 26364 379670 26376
rect 381538 26364 381544 26376
rect 379664 26336 381544 26364
rect 379664 26324 379670 26336
rect 381538 26324 381544 26336
rect 381596 26324 381602 26376
rect 296036 26268 296714 26296
rect 296036 26256 296042 26268
rect 421006 26256 421012 26308
rect 421064 26296 421070 26308
rect 424042 26296 424048 26308
rect 421064 26268 424048 26296
rect 421064 26256 421070 26268
rect 424042 26256 424048 26268
rect 424100 26256 424106 26308
rect 467834 26256 467840 26308
rect 467892 26296 467898 26308
rect 471330 26296 471336 26308
rect 467892 26268 471336 26296
rect 467892 26256 467898 26268
rect 471330 26256 471336 26268
rect 471388 26256 471394 26308
rect 478690 26256 478696 26308
rect 478748 26296 478754 26308
rect 482278 26296 482284 26308
rect 478748 26268 482284 26296
rect 478748 26256 478754 26268
rect 482278 26256 482284 26268
rect 482336 26256 482342 26308
rect 382274 26188 382280 26240
rect 382332 26228 382338 26240
rect 383194 26228 383200 26240
rect 382332 26200 383200 26228
rect 382332 26188 382338 26200
rect 383194 26188 383200 26200
rect 383252 26188 383258 26240
rect 386414 26188 386420 26240
rect 386472 26228 386478 26240
rect 387702 26228 387708 26240
rect 386472 26200 387708 26228
rect 386472 26188 386478 26200
rect 387702 26188 387708 26200
rect 387760 26188 387766 26240
rect 353386 26120 353392 26172
rect 353444 26160 353450 26172
rect 396074 26160 396080 26172
rect 353444 26132 396080 26160
rect 353444 26120 353450 26132
rect 396074 26120 396080 26132
rect 396132 26120 396138 26172
rect 70394 26052 70400 26104
rect 70452 26092 70458 26104
rect 71222 26092 71228 26104
rect 70452 26064 71228 26092
rect 70452 26052 70458 26064
rect 71222 26052 71228 26064
rect 71280 26052 71286 26104
rect 74626 26052 74632 26104
rect 74684 26092 74690 26104
rect 75822 26092 75828 26104
rect 74684 26064 75828 26092
rect 74684 26052 74690 26064
rect 75822 26052 75828 26064
rect 75880 26052 75886 26104
rect 376018 26052 376024 26104
rect 376076 26092 376082 26104
rect 441614 26092 441620 26104
rect 376076 26064 441620 26092
rect 376076 26052 376082 26064
rect 441614 26052 441620 26064
rect 441672 26052 441678 26104
rect 200206 25984 200212 26036
rect 200264 26024 200270 26036
rect 316126 26024 316132 26036
rect 200264 25996 316132 26024
rect 200264 25984 200270 25996
rect 316126 25984 316132 25996
rect 316184 25984 316190 26036
rect 343634 25984 343640 26036
rect 343692 26024 343698 26036
rect 423674 26024 423680 26036
rect 343692 25996 423680 26024
rect 343692 25984 343698 25996
rect 423674 25984 423680 25996
rect 423732 25984 423738 26036
rect 197354 25916 197360 25968
rect 197412 25956 197418 25968
rect 285766 25956 285772 25968
rect 197412 25928 285772 25956
rect 197412 25916 197418 25928
rect 285766 25916 285772 25928
rect 285824 25916 285830 25968
rect 312538 25916 312544 25968
rect 312596 25956 312602 25968
rect 429194 25956 429200 25968
rect 312596 25928 429200 25956
rect 312596 25916 312602 25928
rect 429194 25916 429200 25928
rect 429252 25916 429258 25968
rect 208486 25848 208492 25900
rect 208544 25888 208550 25900
rect 351914 25888 351920 25900
rect 208544 25860 351920 25888
rect 208544 25848 208550 25860
rect 351914 25848 351920 25860
rect 351972 25848 351978 25900
rect 356054 25848 356060 25900
rect 356112 25888 356118 25900
rect 464338 25888 464344 25900
rect 356112 25860 464344 25888
rect 356112 25848 356118 25860
rect 464338 25848 464344 25860
rect 464396 25848 464402 25900
rect 216766 25780 216772 25832
rect 216824 25820 216830 25832
rect 383654 25820 383660 25832
rect 216824 25792 383660 25820
rect 216824 25780 216830 25792
rect 383654 25780 383660 25792
rect 383712 25780 383718 25832
rect 231946 25712 231952 25764
rect 232004 25752 232010 25764
rect 440326 25752 440332 25764
rect 232004 25724 440332 25752
rect 232004 25712 232010 25724
rect 440326 25712 440332 25724
rect 440384 25712 440390 25764
rect 84194 25644 84200 25696
rect 84252 25684 84258 25696
rect 118786 25684 118792 25696
rect 84252 25656 118792 25684
rect 84252 25644 84258 25656
rect 118786 25644 118792 25656
rect 118844 25644 118850 25696
rect 247034 25644 247040 25696
rect 247092 25684 247098 25696
rect 501046 25684 501052 25696
rect 247092 25656 501052 25684
rect 247092 25644 247098 25656
rect 501046 25644 501052 25656
rect 501104 25644 501110 25696
rect 4798 25576 4804 25628
rect 4856 25616 4862 25628
rect 55306 25616 55312 25628
rect 4856 25588 55312 25616
rect 4856 25576 4862 25588
rect 55306 25576 55312 25588
rect 55364 25576 55370 25628
rect 88334 25576 88340 25628
rect 88392 25616 88398 25628
rect 135254 25616 135260 25628
rect 88392 25588 135260 25616
rect 88392 25576 88398 25588
rect 135254 25576 135260 25588
rect 135312 25576 135318 25628
rect 259546 25576 259552 25628
rect 259604 25616 259610 25628
rect 547874 25616 547880 25628
rect 259604 25588 547880 25616
rect 259604 25576 259610 25588
rect 547874 25576 547880 25588
rect 547932 25576 547938 25628
rect 27614 25508 27620 25560
rect 27672 25548 27678 25560
rect 91002 25548 91008 25560
rect 27672 25520 91008 25548
rect 27672 25508 27678 25520
rect 91002 25508 91008 25520
rect 91060 25508 91066 25560
rect 183554 25508 183560 25560
rect 183612 25548 183618 25560
rect 252554 25548 252560 25560
rect 183612 25520 252560 25548
rect 183612 25508 183618 25520
rect 252554 25508 252560 25520
rect 252612 25508 252618 25560
rect 266354 25508 266360 25560
rect 266412 25548 266418 25560
rect 575474 25548 575480 25560
rect 266412 25520 575480 25548
rect 266412 25508 266418 25520
rect 575474 25508 575480 25520
rect 575532 25508 575538 25560
rect 345106 24692 345112 24744
rect 345164 24732 345170 24744
rect 432138 24732 432144 24744
rect 345164 24704 432144 24732
rect 345164 24692 345170 24704
rect 432138 24692 432144 24704
rect 432196 24692 432202 24744
rect 189074 24624 189080 24676
rect 189132 24664 189138 24676
rect 277394 24664 277400 24676
rect 189132 24636 277400 24664
rect 189132 24624 189138 24636
rect 277394 24624 277400 24636
rect 277452 24624 277458 24676
rect 339126 24624 339132 24676
rect 339184 24664 339190 24676
rect 390646 24664 390652 24676
rect 339184 24636 390652 24664
rect 339184 24624 339190 24636
rect 390646 24624 390652 24636
rect 390704 24624 390710 24676
rect 198734 24556 198740 24608
rect 198792 24596 198798 24608
rect 313274 24596 313280 24608
rect 198792 24568 313280 24596
rect 198792 24556 198798 24568
rect 313274 24556 313280 24568
rect 313332 24556 313338 24608
rect 330478 24556 330484 24608
rect 330536 24596 330542 24608
rect 431954 24596 431960 24608
rect 330536 24568 431960 24596
rect 330536 24556 330542 24568
rect 431954 24556 431960 24568
rect 432012 24556 432018 24608
rect 276658 24488 276664 24540
rect 276716 24528 276722 24540
rect 419626 24528 419632 24540
rect 276716 24500 419632 24528
rect 276716 24488 276722 24500
rect 419626 24488 419632 24500
rect 419684 24488 419690 24540
rect 205726 24420 205732 24472
rect 205784 24460 205790 24472
rect 338114 24460 338120 24472
rect 205784 24432 338120 24460
rect 205784 24420 205790 24432
rect 338114 24420 338120 24432
rect 338172 24420 338178 24472
rect 367094 24420 367100 24472
rect 367152 24460 367158 24472
rect 516134 24460 516140 24472
rect 367152 24432 516140 24460
rect 367152 24420 367158 24432
rect 516134 24420 516140 24432
rect 516192 24420 516198 24472
rect 213914 24352 213920 24404
rect 213972 24392 213978 24404
rect 369854 24392 369860 24404
rect 213972 24364 369860 24392
rect 213972 24352 213978 24364
rect 369854 24352 369860 24364
rect 369912 24352 369918 24404
rect 385678 24352 385684 24404
rect 385736 24392 385742 24404
rect 447134 24392 447140 24404
rect 385736 24364 447140 24392
rect 385736 24352 385742 24364
rect 447134 24352 447140 24364
rect 447192 24352 447198 24404
rect 224954 24284 224960 24336
rect 225012 24324 225018 24336
rect 412634 24324 412640 24336
rect 225012 24296 412640 24324
rect 225012 24284 225018 24296
rect 412634 24284 412640 24296
rect 412692 24284 412698 24336
rect 46934 24216 46940 24268
rect 46992 24256 46998 24268
rect 66254 24256 66260 24268
rect 46992 24228 66260 24256
rect 46992 24216 46998 24228
rect 66254 24216 66260 24228
rect 66312 24216 66318 24268
rect 69106 24216 69112 24268
rect 69164 24256 69170 24268
rect 102226 24256 102232 24268
rect 69164 24228 102232 24256
rect 69164 24216 69170 24228
rect 102226 24216 102232 24228
rect 102284 24216 102290 24268
rect 235994 24216 236000 24268
rect 236052 24256 236058 24268
rect 458266 24256 458272 24268
rect 236052 24228 458272 24256
rect 236052 24216 236058 24228
rect 458266 24216 458272 24228
rect 458324 24216 458330 24268
rect 44174 24148 44180 24200
rect 44232 24188 44238 24200
rect 95142 24188 95148 24200
rect 44232 24160 95148 24188
rect 44232 24148 44238 24160
rect 95142 24148 95148 24160
rect 95200 24148 95206 24200
rect 99374 24148 99380 24200
rect 99432 24188 99438 24200
rect 138014 24188 138020 24200
rect 99432 24160 138020 24188
rect 99432 24148 99438 24160
rect 138014 24148 138020 24160
rect 138072 24148 138078 24200
rect 248414 24148 248420 24200
rect 248472 24188 248478 24200
rect 505094 24188 505100 24200
rect 248472 24160 505100 24188
rect 248472 24148 248478 24160
rect 505094 24148 505100 24160
rect 505152 24148 505158 24200
rect 13814 24080 13820 24132
rect 13872 24120 13878 24132
rect 117222 24120 117228 24132
rect 13872 24092 117228 24120
rect 13872 24080 13878 24092
rect 117222 24080 117228 24092
rect 117280 24080 117286 24132
rect 176746 24080 176752 24132
rect 176804 24120 176810 24132
rect 227714 24120 227720 24132
rect 176804 24092 227720 24120
rect 176804 24080 176810 24092
rect 227714 24080 227720 24092
rect 227772 24080 227778 24132
rect 259454 24080 259460 24132
rect 259512 24120 259518 24132
rect 550634 24120 550640 24132
rect 259512 24092 550640 24120
rect 259512 24080 259518 24092
rect 550634 24080 550640 24092
rect 550692 24080 550698 24132
rect 336734 23332 336740 23384
rect 336792 23372 336798 23384
rect 398834 23372 398840 23384
rect 336792 23344 398840 23372
rect 336792 23332 336798 23344
rect 398834 23332 398840 23344
rect 398892 23332 398898 23384
rect 197538 23264 197544 23316
rect 197596 23304 197602 23316
rect 306466 23304 306472 23316
rect 197596 23276 306472 23304
rect 197596 23264 197602 23276
rect 306466 23264 306472 23276
rect 306524 23264 306530 23316
rect 341518 23264 341524 23316
rect 341576 23304 341582 23316
rect 434806 23304 434812 23316
rect 341576 23276 434812 23304
rect 341576 23264 341582 23276
rect 434806 23264 434812 23276
rect 434864 23264 434870 23316
rect 205634 23196 205640 23248
rect 205692 23236 205698 23248
rect 340874 23236 340880 23248
rect 205692 23208 340880 23236
rect 205692 23196 205698 23208
rect 340874 23196 340880 23208
rect 340932 23196 340938 23248
rect 354674 23196 354680 23248
rect 354732 23236 354738 23248
rect 466454 23236 466460 23248
rect 354732 23208 466460 23236
rect 354732 23196 354738 23208
rect 466454 23196 466460 23208
rect 466512 23196 466518 23248
rect 147858 23128 147864 23180
rect 147916 23168 147922 23180
rect 271966 23168 271972 23180
rect 147916 23140 271972 23168
rect 147916 23128 147922 23140
rect 271966 23128 271972 23140
rect 272024 23128 272030 23180
rect 273254 23128 273260 23180
rect 273312 23168 273318 23180
rect 416682 23168 416688 23180
rect 273312 23140 416688 23168
rect 273312 23128 273318 23140
rect 416682 23128 416688 23140
rect 416740 23128 416746 23180
rect 215294 23060 215300 23112
rect 215352 23100 215358 23112
rect 376754 23100 376760 23112
rect 215352 23072 376760 23100
rect 215352 23060 215358 23072
rect 376754 23060 376760 23072
rect 376812 23060 376818 23112
rect 129826 22992 129832 23044
rect 129884 23032 129890 23044
rect 267826 23032 267832 23044
rect 129884 23004 267832 23032
rect 129884 22992 129890 23004
rect 267826 22992 267832 23004
rect 267884 22992 267890 23044
rect 371326 22992 371332 23044
rect 371384 23032 371390 23044
rect 534074 23032 534080 23044
rect 371384 23004 534080 23032
rect 371384 22992 371390 23004
rect 534074 22992 534080 23004
rect 534132 22992 534138 23044
rect 51074 22924 51080 22976
rect 51132 22964 51138 22976
rect 67726 22964 67732 22976
rect 51132 22936 67732 22964
rect 51132 22924 51138 22936
rect 67726 22924 67732 22936
rect 67784 22924 67790 22976
rect 227898 22924 227904 22976
rect 227956 22964 227962 22976
rect 426434 22964 426440 22976
rect 227956 22936 426440 22964
rect 227956 22924 227962 22936
rect 426434 22924 426440 22936
rect 426492 22924 426498 22976
rect 87046 22856 87052 22908
rect 87104 22896 87110 22908
rect 106274 22896 106280 22908
rect 87104 22868 106280 22896
rect 87104 22856 87110 22868
rect 106274 22856 106280 22868
rect 106332 22856 106338 22908
rect 245746 22856 245752 22908
rect 245804 22896 245810 22908
rect 498286 22896 498292 22908
rect 245804 22868 498292 22896
rect 245804 22856 245810 22868
rect 498286 22856 498292 22868
rect 498344 22856 498350 22908
rect 67726 22788 67732 22840
rect 67784 22828 67790 22840
rect 129734 22828 129740 22840
rect 67784 22800 129740 22828
rect 67784 22788 67790 22800
rect 129734 22788 129740 22800
rect 129792 22788 129798 22840
rect 253934 22788 253940 22840
rect 253992 22828 253998 22840
rect 529934 22828 529940 22840
rect 253992 22800 529940 22828
rect 253992 22788 253998 22800
rect 529934 22788 529940 22800
rect 529992 22788 529998 22840
rect 22094 22720 22100 22772
rect 22152 22760 22158 22772
rect 89714 22760 89720 22772
rect 22152 22732 89720 22760
rect 22152 22720 22158 22732
rect 89714 22720 89720 22732
rect 89772 22720 89778 22772
rect 173986 22720 173992 22772
rect 174044 22760 174050 22772
rect 218054 22760 218060 22772
rect 174044 22732 218060 22760
rect 174044 22720 174050 22732
rect 218054 22720 218060 22732
rect 218112 22720 218118 22772
rect 264974 22720 264980 22772
rect 265032 22760 265038 22772
rect 572714 22760 572720 22772
rect 265032 22732 572720 22760
rect 265032 22720 265038 22732
rect 572714 22720 572720 22732
rect 572772 22720 572778 22772
rect 193306 21972 193312 22024
rect 193364 22012 193370 22024
rect 284294 22012 284300 22024
rect 193364 21984 284300 22012
rect 193364 21972 193370 21984
rect 284294 21972 284300 21984
rect 284352 21972 284358 22024
rect 367830 21972 367836 22024
rect 367888 22012 367894 22024
rect 440418 22012 440424 22024
rect 367888 21984 440424 22012
rect 367888 21972 367894 21984
rect 440418 21972 440424 21984
rect 440476 21972 440482 22024
rect 197446 21904 197452 21956
rect 197504 21944 197510 21956
rect 309318 21944 309324 21956
rect 197504 21916 309324 21944
rect 197504 21904 197510 21916
rect 309318 21904 309324 21916
rect 309376 21904 309382 21956
rect 342346 21904 342352 21956
rect 342404 21944 342410 21956
rect 420914 21944 420920 21956
rect 342404 21916 420920 21944
rect 342404 21904 342410 21916
rect 420914 21904 420920 21916
rect 420972 21904 420978 21956
rect 143718 21836 143724 21888
rect 143776 21876 143782 21888
rect 271874 21876 271880 21888
rect 143776 21848 271880 21876
rect 143776 21836 143782 21848
rect 271874 21836 271880 21848
rect 271932 21836 271938 21888
rect 322198 21836 322204 21888
rect 322256 21876 322262 21888
rect 430574 21876 430580 21888
rect 322256 21848 430580 21876
rect 322256 21836 322262 21848
rect 430574 21836 430580 21848
rect 430632 21836 430638 21888
rect 251174 21768 251180 21820
rect 251232 21808 251238 21820
rect 410426 21808 410432 21820
rect 251232 21780 410432 21808
rect 251232 21768 251238 21780
rect 410426 21768 410432 21780
rect 410484 21768 410490 21820
rect 216674 21700 216680 21752
rect 216732 21740 216738 21752
rect 380986 21740 380992 21752
rect 216732 21712 380992 21740
rect 216732 21700 216738 21712
rect 380986 21700 380992 21712
rect 381044 21700 381050 21752
rect 208394 21632 208400 21684
rect 208452 21672 208458 21684
rect 349154 21672 349160 21684
rect 208452 21644 349160 21672
rect 208452 21632 208458 21644
rect 349154 21632 349160 21644
rect 349212 21632 349218 21684
rect 372614 21632 372620 21684
rect 372672 21672 372678 21684
rect 538214 21672 538220 21684
rect 372672 21644 538220 21672
rect 372672 21632 372678 21644
rect 538214 21632 538220 21644
rect 538272 21632 538278 21684
rect 229094 21564 229100 21616
rect 229152 21604 229158 21616
rect 430574 21604 430580 21616
rect 229152 21576 430580 21604
rect 229152 21564 229158 21576
rect 430574 21564 430580 21576
rect 430632 21564 430638 21616
rect 80146 21496 80152 21548
rect 80204 21536 80210 21548
rect 104986 21536 104992 21548
rect 80204 21508 104992 21536
rect 80204 21496 80210 21508
rect 104986 21496 104992 21508
rect 105044 21496 105050 21548
rect 244274 21496 244280 21548
rect 244332 21536 244338 21548
rect 490006 21536 490012 21548
rect 244332 21508 490012 21536
rect 244332 21496 244338 21508
rect 490006 21496 490012 21508
rect 490064 21496 490070 21548
rect 16574 21428 16580 21480
rect 16632 21468 16638 21480
rect 59262 21468 59268 21480
rect 16632 21440 59268 21468
rect 16632 21428 16638 21440
rect 59262 21428 59268 21440
rect 59320 21428 59326 21480
rect 74718 21428 74724 21480
rect 74776 21468 74782 21480
rect 131206 21468 131212 21480
rect 74776 21440 131212 21468
rect 74776 21428 74782 21440
rect 131206 21428 131212 21440
rect 131264 21428 131270 21480
rect 252646 21428 252652 21480
rect 252704 21468 252710 21480
rect 523034 21468 523040 21480
rect 252704 21440 523040 21468
rect 252704 21428 252710 21440
rect 523034 21428 523040 21440
rect 523092 21428 523098 21480
rect 34514 21360 34520 21412
rect 34572 21400 34578 21412
rect 92474 21400 92480 21412
rect 34572 21372 92480 21400
rect 34572 21360 34578 21372
rect 92474 21360 92480 21372
rect 92532 21360 92538 21412
rect 173894 21360 173900 21412
rect 173952 21400 173958 21412
rect 213914 21400 213920 21412
rect 173952 21372 213920 21400
rect 173952 21360 173958 21372
rect 213914 21360 213920 21372
rect 213972 21360 213978 21412
rect 263594 21360 263600 21412
rect 263652 21400 263658 21412
rect 564526 21400 564532 21412
rect 263652 21372 564532 21400
rect 263652 21360 263658 21372
rect 564526 21360 564532 21372
rect 564584 21360 564590 21412
rect 360470 20544 360476 20596
rect 360528 20584 360534 20596
rect 414198 20584 414204 20596
rect 360528 20556 414204 20584
rect 360528 20544 360534 20556
rect 414198 20544 414204 20556
rect 414256 20544 414262 20596
rect 325694 20476 325700 20528
rect 325752 20516 325758 20528
rect 424410 20516 424416 20528
rect 325752 20488 424416 20516
rect 325752 20476 325758 20488
rect 424410 20476 424416 20488
rect 424468 20476 424474 20528
rect 205542 20408 205548 20460
rect 205600 20448 205606 20460
rect 331398 20448 331404 20460
rect 205600 20420 331404 20448
rect 205600 20408 205606 20420
rect 331398 20408 331404 20420
rect 331456 20408 331462 20460
rect 346486 20408 346492 20460
rect 346544 20448 346550 20460
rect 434714 20448 434720 20460
rect 346544 20420 434720 20448
rect 346544 20408 346550 20420
rect 434714 20408 434720 20420
rect 434772 20408 434778 20460
rect 136818 20340 136824 20392
rect 136876 20380 136882 20392
rect 269206 20380 269212 20392
rect 136876 20352 269212 20380
rect 136876 20340 136882 20352
rect 269206 20340 269212 20352
rect 269264 20340 269270 20392
rect 284294 20340 284300 20392
rect 284352 20380 284358 20392
rect 421006 20380 421012 20392
rect 284352 20352 421012 20380
rect 284352 20340 284358 20352
rect 421006 20340 421012 20352
rect 421064 20340 421070 20392
rect 211154 20272 211160 20324
rect 211212 20312 211218 20324
rect 363138 20312 363144 20324
rect 211212 20284 363144 20312
rect 211212 20272 211218 20284
rect 363138 20272 363144 20284
rect 363196 20272 363202 20324
rect 219434 20204 219440 20256
rect 219492 20244 219498 20256
rect 394878 20244 394884 20256
rect 219492 20216 394884 20244
rect 219492 20204 219498 20216
rect 394878 20204 394884 20216
rect 394936 20204 394942 20256
rect 20714 20136 20720 20188
rect 20772 20176 20778 20188
rect 59446 20176 59452 20188
rect 20772 20148 59452 20176
rect 20772 20136 20778 20148
rect 59446 20136 59452 20148
rect 59504 20136 59510 20188
rect 234706 20136 234712 20188
rect 234764 20176 234770 20188
rect 455506 20176 455512 20188
rect 234764 20148 455512 20176
rect 234764 20136 234770 20148
rect 455506 20136 455512 20148
rect 455564 20136 455570 20188
rect 98086 20068 98092 20120
rect 98144 20108 98150 20120
rect 108942 20108 108948 20120
rect 98144 20080 108948 20108
rect 98144 20068 98150 20080
rect 108942 20068 108948 20080
rect 109000 20068 109006 20120
rect 245654 20068 245660 20120
rect 245712 20108 245718 20120
rect 494238 20108 494244 20120
rect 245712 20080 494244 20108
rect 245712 20068 245718 20080
rect 494238 20068 494244 20080
rect 494296 20068 494302 20120
rect 59354 20000 59360 20052
rect 59412 20040 59418 20052
rect 99282 20040 99288 20052
rect 59412 20012 99288 20040
rect 59412 20000 59418 20012
rect 99282 20000 99288 20012
rect 99340 20000 99346 20052
rect 172514 20000 172520 20052
rect 172572 20040 172578 20052
rect 209866 20040 209872 20052
rect 172572 20012 209872 20040
rect 172572 20000 172578 20012
rect 209866 20000 209872 20012
rect 209924 20000 209930 20052
rect 256602 20000 256608 20052
rect 256660 20040 256666 20052
rect 525794 20040 525800 20052
rect 256660 20012 525800 20040
rect 256660 20000 256666 20012
rect 525794 20000 525800 20012
rect 525852 20000 525858 20052
rect 52454 19932 52460 19984
rect 52512 19972 52518 19984
rect 125686 19972 125692 19984
rect 52512 19944 125692 19972
rect 52512 19932 52518 19944
rect 125686 19932 125692 19944
rect 125744 19932 125750 19984
rect 186314 19932 186320 19984
rect 186372 19972 186378 19984
rect 263594 19972 263600 19984
rect 186372 19944 263600 19972
rect 186372 19932 186378 19944
rect 263594 19932 263600 19944
rect 263652 19932 263658 19984
rect 267642 19932 267648 19984
rect 267700 19972 267706 19984
rect 568574 19972 568580 19984
rect 267700 19944 568580 19972
rect 267700 19932 267706 19944
rect 568574 19932 568580 19944
rect 568632 19932 568638 19984
rect 342254 19184 342260 19236
rect 342312 19224 342318 19236
rect 416958 19224 416964 19236
rect 342312 19196 416964 19224
rect 342312 19184 342318 19196
rect 416958 19184 416964 19196
rect 417016 19184 417022 19236
rect 364978 19116 364984 19168
rect 365036 19156 365042 19168
rect 441614 19156 441620 19168
rect 365036 19128 441620 19156
rect 365036 19116 365042 19128
rect 441614 19116 441620 19128
rect 441672 19116 441678 19168
rect 140866 19048 140872 19100
rect 140924 19088 140930 19100
rect 270494 19088 270500 19100
rect 140924 19060 270500 19088
rect 140924 19048 140930 19060
rect 270494 19048 270500 19060
rect 270552 19048 270558 19100
rect 304258 19048 304264 19100
rect 304316 19088 304322 19100
rect 426526 19088 426532 19100
rect 304316 19060 426532 19088
rect 304316 19048 304322 19060
rect 426526 19048 426532 19060
rect 426584 19048 426590 19100
rect 204254 18980 204260 19032
rect 204312 19020 204318 19032
rect 334158 19020 334164 19032
rect 204312 18992 334164 19020
rect 204312 18980 204318 18992
rect 334158 18980 334164 18992
rect 334216 18980 334222 19032
rect 353938 18980 353944 19032
rect 353996 19020 354002 19032
rect 437566 19020 437572 19032
rect 353996 18992 437572 19020
rect 353996 18980 354002 18992
rect 437566 18980 437572 18992
rect 437624 18980 437630 19032
rect 212534 18912 212540 18964
rect 212592 18952 212598 18964
rect 365898 18952 365904 18964
rect 212592 18924 365904 18952
rect 212592 18912 212598 18924
rect 365898 18912 365904 18924
rect 365956 18912 365962 18964
rect 28994 18844 29000 18896
rect 29052 18884 29058 18896
rect 62206 18884 62212 18896
rect 29052 18856 62212 18884
rect 29052 18844 29058 18856
rect 62206 18844 62212 18856
rect 62264 18844 62270 18896
rect 220814 18844 220820 18896
rect 220872 18884 220878 18896
rect 398926 18884 398932 18896
rect 220872 18856 398932 18884
rect 220872 18844 220878 18856
rect 398926 18844 398932 18856
rect 398984 18844 398990 18896
rect 237466 18776 237472 18828
rect 237524 18816 237530 18828
rect 462406 18816 462412 18828
rect 237524 18788 462412 18816
rect 237524 18776 237530 18788
rect 462406 18776 462412 18788
rect 462464 18776 462470 18828
rect 62206 18708 62212 18760
rect 62264 18748 62270 18760
rect 99466 18748 99472 18760
rect 62264 18720 99472 18748
rect 62264 18708 62270 18720
rect 99466 18708 99472 18720
rect 99524 18708 99530 18760
rect 242894 18708 242900 18760
rect 242952 18748 242958 18760
rect 487154 18748 487160 18760
rect 242952 18720 487160 18748
rect 242952 18708 242958 18720
rect 487154 18708 487160 18720
rect 487212 18708 487218 18760
rect 487246 18708 487252 18760
rect 487304 18748 487310 18760
rect 531314 18748 531320 18760
rect 487304 18720 531320 18748
rect 487304 18708 487310 18720
rect 531314 18708 531320 18720
rect 531372 18708 531378 18760
rect 92474 18640 92480 18692
rect 92532 18680 92538 18692
rect 136726 18680 136732 18692
rect 92532 18652 136732 18680
rect 92532 18640 92538 18652
rect 136726 18640 136732 18652
rect 136784 18640 136790 18692
rect 169754 18640 169760 18692
rect 169812 18680 169818 18692
rect 200206 18680 200212 18692
rect 169812 18652 200212 18680
rect 169812 18640 169818 18652
rect 200206 18640 200212 18652
rect 200264 18640 200270 18692
rect 251358 18640 251364 18692
rect 251416 18680 251422 18692
rect 518894 18680 518900 18692
rect 251416 18652 518900 18680
rect 251416 18640 251422 18652
rect 518894 18640 518900 18652
rect 518952 18640 518958 18692
rect 49694 18572 49700 18624
rect 49752 18612 49758 18624
rect 125594 18612 125600 18624
rect 49752 18584 125600 18612
rect 49752 18572 49758 18584
rect 125594 18572 125600 18584
rect 125652 18572 125658 18624
rect 186958 18572 186964 18624
rect 187016 18612 187022 18624
rect 259454 18612 259460 18624
rect 187016 18584 259460 18612
rect 187016 18572 187022 18584
rect 259454 18572 259460 18584
rect 259512 18572 259518 18624
rect 262306 18572 262312 18624
rect 262364 18612 262370 18624
rect 561674 18612 561680 18624
rect 262364 18584 561680 18612
rect 262364 18572 262370 18584
rect 561674 18572 561680 18584
rect 561732 18572 561738 18624
rect 211154 17756 211160 17808
rect 211212 17796 211218 17808
rect 288526 17796 288532 17808
rect 211212 17768 288532 17796
rect 211212 17756 211218 17768
rect 288526 17756 288532 17768
rect 288584 17756 288590 17808
rect 345014 17756 345020 17808
rect 345072 17796 345078 17808
rect 427814 17796 427820 17808
rect 345072 17768 427820 17796
rect 345072 17756 345078 17768
rect 427814 17756 427820 17768
rect 427872 17756 427878 17808
rect 201586 17688 201592 17740
rect 201644 17728 201650 17740
rect 324406 17728 324412 17740
rect 201644 17700 324412 17728
rect 201644 17688 201650 17700
rect 324406 17688 324412 17700
rect 324464 17688 324470 17740
rect 324958 17688 324964 17740
rect 325016 17728 325022 17740
rect 432046 17728 432052 17740
rect 325016 17700 432052 17728
rect 325016 17688 325022 17700
rect 432046 17688 432052 17700
rect 432104 17688 432110 17740
rect 211246 17620 211252 17672
rect 211304 17660 211310 17672
rect 358906 17660 358912 17672
rect 211304 17632 358912 17660
rect 211304 17620 211310 17632
rect 358906 17620 358912 17632
rect 358964 17620 358970 17672
rect 374086 17620 374092 17672
rect 374144 17660 374150 17672
rect 540974 17660 540980 17672
rect 374144 17632 540980 17660
rect 374144 17620 374150 17632
rect 540974 17620 540980 17632
rect 541032 17620 541038 17672
rect 218146 17552 218152 17604
rect 218204 17592 218210 17604
rect 387886 17592 387892 17604
rect 218204 17564 387892 17592
rect 218204 17552 218210 17564
rect 387886 17552 387892 17564
rect 387944 17552 387950 17604
rect 226426 17484 226432 17536
rect 226484 17524 226490 17536
rect 408586 17524 408592 17536
rect 226484 17496 408592 17524
rect 226484 17484 226490 17496
rect 408586 17484 408592 17496
rect 408644 17484 408650 17536
rect 233234 17416 233240 17468
rect 233292 17456 233298 17468
rect 448790 17456 448796 17468
rect 233292 17428 448796 17456
rect 233292 17416 233298 17428
rect 448790 17416 448796 17428
rect 448848 17416 448854 17468
rect 73154 17348 73160 17400
rect 73212 17388 73218 17400
rect 102134 17388 102140 17400
rect 73212 17360 102140 17388
rect 73212 17348 73218 17360
rect 102134 17348 102140 17360
rect 102192 17348 102198 17400
rect 244918 17348 244924 17400
rect 244976 17388 244982 17400
rect 483198 17388 483204 17400
rect 244976 17360 483204 17388
rect 244976 17348 244982 17360
rect 483198 17348 483204 17360
rect 483256 17348 483262 17400
rect 35894 17280 35900 17332
rect 35952 17320 35958 17332
rect 63494 17320 63500 17332
rect 35952 17292 63500 17320
rect 35952 17280 35958 17292
rect 63494 17280 63500 17292
rect 63552 17280 63558 17332
rect 81526 17280 81532 17332
rect 81584 17320 81590 17332
rect 133966 17320 133972 17332
rect 81584 17292 133972 17320
rect 81584 17280 81590 17292
rect 133966 17280 133972 17292
rect 134024 17280 134030 17332
rect 168466 17280 168472 17332
rect 168524 17320 168530 17332
rect 195974 17320 195980 17332
rect 168524 17292 195980 17320
rect 168524 17280 168530 17292
rect 195974 17280 195980 17292
rect 196032 17280 196038 17332
rect 251266 17280 251272 17332
rect 251324 17320 251330 17332
rect 514754 17320 514760 17332
rect 251324 17292 514760 17320
rect 251324 17280 251330 17292
rect 514754 17280 514760 17292
rect 514812 17280 514818 17332
rect 41414 17212 41420 17264
rect 41472 17252 41478 17264
rect 93946 17252 93952 17264
rect 41472 17224 93952 17252
rect 41472 17212 41478 17224
rect 93946 17212 93952 17224
rect 94004 17212 94010 17264
rect 180794 17212 180800 17264
rect 180852 17252 180858 17264
rect 242894 17252 242900 17264
rect 180852 17224 242900 17252
rect 180852 17212 180858 17224
rect 242894 17212 242900 17224
rect 242952 17212 242958 17264
rect 262214 17212 262220 17264
rect 262272 17252 262278 17264
rect 557534 17252 557540 17264
rect 262272 17224 557540 17252
rect 262272 17212 262278 17224
rect 557534 17212 557540 17224
rect 557592 17212 557598 17264
rect 411898 16532 411904 16584
rect 411956 16572 411962 16584
rect 448606 16572 448612 16584
rect 411956 16544 448612 16572
rect 411956 16532 411962 16544
rect 448606 16532 448612 16544
rect 448664 16532 448670 16584
rect 208578 16464 208584 16516
rect 208636 16504 208642 16516
rect 288434 16504 288440 16516
rect 208636 16476 288440 16504
rect 208636 16464 208642 16476
rect 288434 16464 288440 16476
rect 288492 16464 288498 16516
rect 342898 16464 342904 16516
rect 342956 16504 342962 16516
rect 436186 16504 436192 16516
rect 342956 16476 436192 16504
rect 342956 16464 342962 16476
rect 436186 16464 436192 16476
rect 436244 16464 436250 16516
rect 183738 16396 183744 16448
rect 183796 16436 183802 16448
rect 281534 16436 281540 16448
rect 183796 16408 281540 16436
rect 183796 16396 183802 16408
rect 281534 16396 281540 16408
rect 281592 16396 281598 16448
rect 357526 16396 357532 16448
rect 357584 16436 357590 16448
rect 461670 16436 461676 16448
rect 357584 16408 461676 16436
rect 357584 16396 357590 16408
rect 461670 16396 461676 16408
rect 461728 16396 461734 16448
rect 259546 16328 259552 16380
rect 259604 16368 259610 16380
rect 416866 16368 416872 16380
rect 259604 16340 416872 16368
rect 259604 16328 259610 16340
rect 416866 16328 416872 16340
rect 416924 16328 416930 16380
rect 255866 16260 255872 16312
rect 255924 16300 255930 16312
rect 416774 16300 416780 16312
rect 255924 16272 416780 16300
rect 255924 16260 255930 16272
rect 416774 16260 416780 16272
rect 416832 16260 416838 16312
rect 248414 16192 248420 16244
rect 248472 16232 248478 16244
rect 414106 16232 414112 16244
rect 248472 16204 414112 16232
rect 248472 16192 248478 16204
rect 414106 16192 414112 16204
rect 414164 16192 414170 16244
rect 245194 16124 245200 16176
rect 245252 16164 245258 16176
rect 414014 16164 414020 16176
rect 245252 16136 414020 16164
rect 245252 16124 245258 16136
rect 414014 16124 414020 16136
rect 414072 16124 414078 16176
rect 126974 16056 126980 16108
rect 127032 16096 127038 16108
rect 267734 16096 267740 16108
rect 127032 16068 267740 16096
rect 127032 16056 127038 16068
rect 267734 16056 267740 16068
rect 267792 16056 267798 16108
rect 373994 16056 374000 16108
rect 374052 16096 374058 16108
rect 545482 16096 545488 16108
rect 374052 16068 545488 16096
rect 374052 16056 374058 16068
rect 545482 16056 545488 16068
rect 545540 16056 545546 16108
rect 241698 15988 241704 16040
rect 241756 16028 241762 16040
rect 412726 16028 412732 16040
rect 241756 16000 412732 16028
rect 241756 15988 241762 16000
rect 412726 15988 412732 16000
rect 412784 15988 412790 16040
rect 40218 15920 40224 15972
rect 40276 15960 40282 15972
rect 64966 15960 64972 15972
rect 40276 15932 64972 15960
rect 40276 15920 40282 15932
rect 64966 15920 64972 15932
rect 65024 15920 65030 15972
rect 66714 15920 66720 15972
rect 66772 15960 66778 15972
rect 100754 15960 100760 15972
rect 66772 15932 100760 15960
rect 66772 15920 66778 15932
rect 100754 15920 100760 15932
rect 100812 15920 100818 15972
rect 102226 15920 102232 15972
rect 102284 15960 102290 15972
rect 110506 15960 110512 15972
rect 102284 15932 110512 15960
rect 102284 15920 102290 15932
rect 110506 15920 110512 15932
rect 110564 15920 110570 15972
rect 132954 15920 132960 15972
rect 133012 15960 133018 15972
rect 151906 15960 151912 15972
rect 133012 15932 151912 15960
rect 133012 15920 133018 15932
rect 151906 15920 151912 15932
rect 151964 15920 151970 15972
rect 168374 15920 168380 15972
rect 168432 15960 168438 15972
rect 193398 15960 193404 15972
rect 168432 15932 193404 15960
rect 168432 15920 168438 15932
rect 193398 15920 193404 15932
rect 193456 15920 193462 15972
rect 237650 15920 237656 15972
rect 237708 15960 237714 15972
rect 411346 15960 411352 15972
rect 237708 15932 411352 15960
rect 237708 15920 237714 15932
rect 411346 15920 411352 15932
rect 411404 15920 411410 15972
rect 418890 15920 418896 15972
rect 418948 15960 418954 15972
rect 473446 15960 473452 15972
rect 418948 15932 473452 15960
rect 418948 15920 418954 15932
rect 473446 15920 473452 15932
rect 473504 15920 473510 15972
rect 488626 15920 488632 15972
rect 488684 15960 488690 15972
rect 536098 15960 536104 15972
rect 488684 15932 536104 15960
rect 488684 15920 488690 15932
rect 536098 15920 536104 15932
rect 536156 15920 536162 15972
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 116026 15892 116032 15904
rect 11756 15864 116032 15892
rect 11756 15852 11762 15864
rect 116026 15852 116032 15864
rect 116084 15852 116090 15904
rect 138842 15852 138848 15904
rect 138900 15892 138906 15904
rect 386506 15892 386512 15904
rect 138900 15864 386512 15892
rect 138900 15852 138906 15864
rect 386506 15852 386512 15864
rect 386564 15852 386570 15904
rect 414658 15852 414664 15904
rect 414716 15892 414722 15904
rect 520274 15892 520280 15904
rect 414716 15864 520280 15892
rect 414716 15852 414722 15864
rect 520274 15852 520280 15864
rect 520332 15852 520338 15904
rect 378778 15104 378784 15156
rect 378836 15144 378842 15156
rect 443086 15144 443092 15156
rect 378836 15116 443092 15144
rect 378836 15104 378842 15116
rect 443086 15104 443092 15116
rect 443144 15104 443150 15156
rect 335998 15036 336004 15088
rect 336056 15076 336062 15088
rect 433334 15076 433340 15088
rect 336056 15048 433340 15076
rect 336056 15036 336062 15048
rect 433334 15036 433340 15048
rect 433392 15036 433398 15088
rect 294598 14968 294604 15020
rect 294656 15008 294662 15020
rect 425146 15008 425152 15020
rect 294656 14980 425152 15008
rect 294656 14968 294662 14980
rect 425146 14968 425152 14980
rect 425204 14968 425210 15020
rect 231026 14900 231032 14952
rect 231084 14940 231090 14952
rect 409874 14940 409880 14952
rect 231084 14912 409880 14940
rect 231084 14900 231090 14912
rect 409874 14900 409880 14912
rect 409932 14900 409938 14952
rect 381538 14832 381544 14884
rect 381596 14872 381602 14884
rect 563054 14872 563060 14884
rect 381596 14844 563060 14872
rect 381596 14832 381602 14844
rect 563054 14832 563060 14844
rect 563112 14832 563118 14884
rect 219986 14764 219992 14816
rect 220044 14804 220050 14816
rect 407114 14804 407120 14816
rect 220044 14776 407120 14804
rect 220044 14764 220050 14776
rect 407114 14764 407120 14776
rect 407172 14764 407178 14816
rect 216858 14696 216864 14748
rect 216916 14736 216922 14748
rect 405734 14736 405740 14748
rect 216916 14708 405740 14736
rect 216916 14696 216922 14708
rect 405734 14696 405740 14708
rect 405792 14696 405798 14748
rect 213362 14628 213368 14680
rect 213420 14668 213426 14680
rect 405826 14668 405832 14680
rect 213420 14640 405832 14668
rect 213420 14628 213426 14640
rect 405826 14628 405832 14640
rect 405884 14628 405890 14680
rect 82906 14560 82912 14612
rect 82964 14600 82970 14612
rect 111610 14600 111616 14612
rect 82964 14572 111616 14600
rect 82964 14560 82970 14572
rect 111610 14560 111616 14572
rect 111668 14560 111674 14612
rect 209958 14560 209964 14612
rect 210016 14600 210022 14612
rect 404354 14600 404360 14612
rect 210016 14572 404360 14600
rect 210016 14560 210022 14572
rect 404354 14560 404360 14572
rect 404412 14560 404418 14612
rect 404998 14560 405004 14612
rect 405056 14600 405062 14612
rect 445846 14600 445852 14612
rect 405056 14572 445852 14600
rect 405056 14560 405062 14572
rect 445846 14560 445852 14572
rect 445904 14560 445910 14612
rect 60826 14492 60832 14544
rect 60884 14532 60890 14544
rect 128446 14532 128452 14544
rect 60884 14504 128452 14532
rect 60884 14492 60890 14504
rect 128446 14492 128452 14504
rect 128504 14492 128510 14544
rect 206186 14492 206192 14544
rect 206244 14532 206250 14544
rect 403066 14532 403072 14544
rect 206244 14504 403072 14532
rect 206244 14492 206250 14504
rect 403066 14492 403072 14504
rect 403124 14492 403130 14544
rect 410518 14492 410524 14544
rect 410576 14532 410582 14544
rect 495526 14532 495532 14544
rect 410576 14504 495532 14532
rect 410576 14492 410582 14504
rect 495526 14492 495532 14504
rect 495584 14492 495590 14544
rect 14458 14424 14464 14476
rect 14516 14464 14522 14476
rect 88518 14464 88524 14476
rect 14516 14436 88524 14464
rect 14516 14424 14522 14436
rect 88518 14424 88524 14436
rect 88576 14424 88582 14476
rect 135254 14424 135260 14476
rect 135312 14464 135318 14476
rect 385126 14464 385132 14476
rect 135312 14436 385132 14464
rect 135312 14424 135318 14436
rect 385126 14424 385132 14436
rect 385184 14424 385190 14476
rect 407850 14424 407856 14476
rect 407908 14464 407914 14476
rect 554774 14464 554780 14476
rect 407908 14436 554780 14464
rect 407908 14424 407914 14436
rect 554774 14424 554780 14436
rect 554832 14424 554838 14476
rect 268378 13676 268384 13728
rect 268436 13716 268442 13728
rect 303614 13716 303620 13728
rect 268436 13688 303620 13716
rect 268436 13676 268442 13688
rect 303614 13676 303620 13688
rect 303672 13676 303678 13728
rect 346394 13676 346400 13728
rect 346452 13716 346458 13728
rect 439130 13716 439136 13728
rect 346452 13688 439136 13716
rect 346452 13676 346458 13688
rect 439130 13676 439136 13688
rect 439188 13676 439194 13728
rect 273898 13608 273904 13660
rect 273956 13648 273962 13660
rect 374086 13648 374092 13660
rect 273956 13620 374092 13648
rect 273956 13608 273962 13620
rect 374086 13608 374092 13620
rect 374144 13608 374150 13660
rect 158898 13540 158904 13592
rect 158956 13580 158962 13592
rect 274634 13580 274640 13592
rect 158956 13552 274640 13580
rect 158956 13540 158962 13552
rect 274634 13540 274640 13552
rect 274692 13540 274698 13592
rect 376110 13540 376116 13592
rect 376168 13580 376174 13592
rect 492306 13580 492312 13592
rect 376168 13552 492312 13580
rect 376168 13540 376174 13552
rect 492306 13540 492312 13552
rect 492364 13540 492370 13592
rect 154666 13472 154672 13524
rect 154724 13512 154730 13524
rect 274726 13512 274732 13524
rect 154724 13484 274732 13512
rect 154724 13472 154730 13484
rect 274726 13472 274732 13484
rect 274784 13472 274790 13524
rect 284938 13472 284944 13524
rect 284996 13512 285002 13524
rect 422386 13512 422392 13524
rect 284996 13484 422392 13512
rect 284996 13472 285002 13484
rect 422386 13472 422392 13484
rect 422444 13472 422450 13524
rect 151998 13404 152004 13456
rect 152056 13444 152062 13456
rect 273346 13444 273352 13456
rect 152056 13416 273352 13444
rect 152056 13404 152062 13416
rect 273346 13404 273352 13416
rect 273404 13404 273410 13456
rect 369946 13404 369952 13456
rect 370004 13444 370010 13456
rect 527818 13444 527824 13456
rect 370004 13416 527824 13444
rect 370004 13404 370010 13416
rect 527818 13404 527824 13416
rect 527876 13404 527882 13456
rect 249058 13336 249064 13388
rect 249116 13376 249122 13388
rect 415394 13376 415400 13388
rect 249116 13348 415400 13376
rect 249116 13336 249122 13348
rect 415394 13336 415400 13348
rect 415452 13336 415458 13388
rect 234614 13268 234620 13320
rect 234672 13308 234678 13320
rect 451642 13308 451648 13320
rect 234672 13280 451648 13308
rect 234672 13268 234678 13280
rect 451642 13268 451648 13280
rect 451700 13268 451706 13320
rect 80238 13200 80244 13252
rect 80296 13240 80302 13252
rect 100754 13240 100760 13252
rect 80296 13212 100760 13240
rect 80296 13200 80302 13212
rect 100754 13200 100760 13212
rect 100812 13200 100818 13252
rect 173894 13200 173900 13252
rect 173952 13240 173958 13252
rect 394786 13240 394792 13252
rect 173952 13212 394792 13240
rect 173952 13200 173958 13212
rect 394786 13200 394792 13212
rect 394844 13200 394850 13252
rect 64322 13132 64328 13184
rect 64380 13172 64386 13184
rect 128354 13172 128360 13184
rect 64380 13144 128360 13172
rect 64380 13132 64386 13144
rect 128354 13132 128360 13144
rect 128412 13132 128418 13184
rect 170306 13132 170312 13184
rect 170364 13172 170370 13184
rect 394694 13172 394700 13184
rect 170364 13144 394700 13172
rect 170364 13132 170370 13144
rect 394694 13132 394700 13144
rect 394752 13132 394758 13184
rect 485774 13132 485780 13184
rect 485832 13172 485838 13184
rect 528554 13172 528560 13184
rect 485832 13144 528560 13172
rect 485832 13132 485838 13144
rect 528554 13132 528560 13144
rect 528612 13132 528618 13184
rect 17954 13064 17960 13116
rect 18012 13104 18018 13116
rect 88426 13104 88432 13116
rect 18012 13076 88432 13104
rect 18012 13064 18018 13076
rect 88426 13064 88432 13076
rect 88484 13064 88490 13116
rect 128170 13064 128176 13116
rect 128228 13104 128234 13116
rect 383746 13104 383752 13116
rect 128228 13076 383752 13104
rect 128228 13064 128234 13076
rect 383746 13064 383752 13076
rect 383804 13064 383810 13116
rect 396810 13064 396816 13116
rect 396868 13104 396874 13116
rect 508866 13104 508872 13116
rect 396868 13076 508872 13104
rect 396868 13064 396874 13076
rect 508866 13064 508872 13076
rect 508924 13064 508930 13116
rect 360838 12996 360844 13048
rect 360896 13036 360902 13048
rect 438854 13036 438860 13048
rect 360896 13008 438860 13036
rect 360896 12996 360902 13008
rect 438854 12996 438860 13008
rect 438912 12996 438918 13048
rect 105722 12452 105728 12504
rect 105780 12492 105786 12504
rect 110414 12492 110420 12504
rect 105780 12464 110420 12492
rect 105780 12452 105786 12464
rect 110414 12452 110420 12464
rect 110472 12452 110478 12504
rect 327718 12384 327724 12436
rect 327776 12424 327782 12436
rect 353570 12424 353576 12436
rect 327776 12396 353576 12424
rect 327776 12384 327782 12396
rect 353570 12384 353576 12396
rect 353628 12384 353634 12436
rect 261754 12316 261760 12368
rect 261812 12356 261818 12368
rect 302326 12356 302332 12368
rect 261812 12328 302332 12356
rect 261812 12316 261818 12328
rect 302326 12316 302332 12328
rect 302384 12316 302390 12368
rect 325786 12316 325792 12368
rect 325844 12356 325850 12368
rect 357526 12356 357532 12368
rect 325844 12328 357532 12356
rect 325844 12316 325850 12328
rect 357526 12316 357532 12328
rect 357584 12316 357590 12368
rect 247586 12248 247592 12300
rect 247644 12288 247650 12300
rect 298094 12288 298100 12300
rect 247644 12260 298100 12288
rect 247644 12248 247650 12260
rect 298094 12248 298100 12260
rect 298152 12248 298158 12300
rect 349246 12248 349252 12300
rect 349304 12288 349310 12300
rect 445846 12288 445852 12300
rect 349304 12260 445852 12288
rect 349304 12248 349310 12260
rect 445846 12248 445852 12260
rect 445904 12248 445910 12300
rect 236546 12180 236552 12232
rect 236604 12220 236610 12232
rect 295334 12220 295340 12232
rect 236604 12192 295340 12220
rect 236604 12180 236610 12192
rect 295334 12180 295340 12192
rect 295392 12180 295398 12232
rect 349338 12180 349344 12232
rect 349396 12220 349402 12232
rect 448698 12220 448704 12232
rect 349396 12192 448704 12220
rect 349396 12180 349402 12192
rect 448698 12180 448704 12192
rect 448756 12180 448762 12232
rect 233418 12112 233424 12164
rect 233476 12152 233482 12164
rect 294046 12152 294052 12164
rect 233476 12124 294052 12152
rect 233476 12112 233482 12124
rect 294046 12112 294052 12124
rect 294104 12112 294110 12164
rect 350534 12112 350540 12164
rect 350592 12152 350598 12164
rect 453298 12152 453304 12164
rect 350592 12124 453304 12152
rect 350592 12112 350598 12124
rect 453298 12112 453304 12124
rect 453356 12112 453362 12164
rect 226518 12044 226524 12096
rect 226576 12084 226582 12096
rect 292574 12084 292580 12096
rect 226576 12056 292580 12084
rect 226576 12044 226582 12056
rect 292574 12044 292580 12056
rect 292632 12044 292638 12096
rect 299566 12044 299572 12096
rect 299624 12084 299630 12096
rect 311986 12084 311992 12096
rect 299624 12056 311992 12084
rect 299624 12044 299630 12056
rect 311986 12044 311992 12056
rect 312044 12044 312050 12096
rect 352098 12044 352104 12096
rect 352156 12084 352162 12096
rect 457070 12084 457076 12096
rect 352156 12056 457076 12084
rect 352156 12044 352162 12056
rect 457070 12044 457076 12056
rect 457128 12044 457134 12096
rect 222746 11976 222752 12028
rect 222804 12016 222810 12028
rect 291194 12016 291200 12028
rect 222804 11988 291200 12016
rect 222804 11976 222810 11988
rect 291194 11976 291200 11988
rect 291252 11976 291258 12028
rect 296070 11976 296076 12028
rect 296128 12016 296134 12028
rect 327994 12016 328000 12028
rect 296128 11988 328000 12016
rect 296128 11976 296134 11988
rect 327994 11976 328000 11988
rect 328052 11976 328058 12028
rect 352006 11976 352012 12028
rect 352064 12016 352070 12028
rect 459922 12016 459928 12028
rect 352064 11988 459928 12016
rect 352064 11976 352070 11988
rect 459922 11976 459928 11988
rect 459980 11976 459986 12028
rect 77294 11908 77300 11960
rect 77352 11948 77358 11960
rect 93946 11948 93952 11960
rect 77352 11920 93952 11948
rect 77352 11908 77358 11920
rect 93946 11908 93952 11920
rect 94004 11908 94010 11960
rect 219250 11908 219256 11960
rect 219308 11948 219314 11960
rect 291286 11948 291292 11960
rect 219308 11920 291292 11948
rect 219308 11908 219314 11920
rect 291286 11908 291292 11920
rect 291344 11908 291350 11960
rect 291838 11908 291844 11960
rect 291896 11948 291902 11960
rect 345290 11948 345296 11960
rect 291896 11920 345296 11948
rect 291896 11908 291902 11920
rect 345290 11908 345296 11920
rect 345348 11908 345354 11960
rect 353294 11908 353300 11960
rect 353352 11948 353358 11960
rect 463970 11948 463976 11960
rect 353352 11920 463976 11948
rect 353352 11908 353358 11920
rect 463970 11908 463976 11920
rect 464028 11908 464034 11960
rect 84194 11840 84200 11892
rect 84252 11880 84258 11892
rect 104894 11880 104900 11892
rect 84252 11852 104900 11880
rect 84252 11840 84258 11852
rect 104894 11840 104900 11852
rect 104952 11840 104958 11892
rect 215294 11840 215300 11892
rect 215352 11880 215358 11892
rect 289814 11880 289820 11892
rect 215352 11852 289820 11880
rect 215352 11840 215358 11852
rect 289814 11840 289820 11852
rect 289872 11840 289878 11892
rect 294506 11840 294512 11892
rect 294564 11880 294570 11892
rect 413278 11880 413284 11892
rect 294564 11852 413284 11880
rect 294564 11840 294570 11852
rect 413278 11840 413284 11852
rect 413336 11840 413342 11892
rect 485038 11840 485044 11892
rect 485096 11880 485102 11892
rect 507210 11880 507216 11892
rect 485096 11852 507216 11880
rect 485096 11840 485102 11852
rect 507210 11840 507216 11852
rect 507268 11840 507274 11892
rect 44266 11772 44272 11824
rect 44324 11812 44330 11824
rect 64874 11812 64880 11824
rect 44324 11784 64880 11812
rect 44324 11772 44330 11784
rect 64874 11772 64880 11784
rect 64932 11772 64938 11824
rect 85758 11772 85764 11824
rect 85816 11812 85822 11824
rect 133874 11812 133880 11824
rect 85816 11784 133880 11812
rect 85816 11772 85822 11784
rect 133874 11772 133880 11784
rect 133932 11772 133938 11824
rect 133966 11772 133972 11824
rect 134024 11812 134030 11824
rect 269114 11812 269120 11824
rect 134024 11784 269120 11812
rect 134024 11772 134030 11784
rect 269114 11772 269120 11784
rect 269172 11772 269178 11824
rect 273898 11772 273904 11824
rect 273956 11812 273962 11824
rect 418154 11812 418160 11824
rect 273956 11784 418160 11812
rect 273956 11772 273962 11784
rect 418154 11772 418160 11784
rect 418212 11772 418218 11824
rect 484394 11772 484400 11824
rect 484452 11812 484458 11824
rect 521654 11812 521660 11824
rect 484452 11784 521660 11812
rect 484452 11772 484458 11784
rect 521654 11772 521660 11784
rect 521712 11772 521718 11824
rect 30834 11704 30840 11756
rect 30892 11744 30898 11756
rect 90358 11744 90364 11756
rect 30892 11716 90364 11744
rect 30892 11704 30898 11716
rect 90358 11704 90364 11716
rect 90416 11704 90422 11756
rect 188522 11704 188528 11756
rect 188580 11744 188586 11756
rect 399018 11744 399024 11756
rect 188580 11716 399024 11744
rect 188580 11704 188586 11716
rect 399018 11704 399024 11716
rect 399076 11704 399082 11756
rect 453390 11704 453396 11756
rect 453448 11744 453454 11756
rect 566826 11744 566832 11756
rect 453448 11716 566832 11744
rect 453448 11704 453454 11716
rect 566826 11704 566832 11716
rect 566884 11704 566890 11756
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 264974 10956 264980 11008
rect 265032 10996 265038 11008
rect 302234 10996 302240 11008
rect 265032 10968 302240 10996
rect 265032 10956 265038 10968
rect 302234 10956 302240 10968
rect 302292 10956 302298 11008
rect 311434 10956 311440 11008
rect 311492 10996 311498 11008
rect 313918 10996 313924 11008
rect 311492 10968 313924 10996
rect 311492 10956 311498 10968
rect 313918 10956 313924 10968
rect 313976 10956 313982 11008
rect 334066 10956 334072 11008
rect 334124 10996 334130 11008
rect 389450 10996 389456 11008
rect 334124 10968 389456 10996
rect 334124 10956 334130 10968
rect 389450 10956 389456 10968
rect 389508 10956 389514 11008
rect 251266 10888 251272 10940
rect 251324 10928 251330 10940
rect 299658 10928 299664 10940
rect 251324 10900 299664 10928
rect 251324 10888 251330 10900
rect 299658 10888 299664 10900
rect 299716 10888 299722 10940
rect 335354 10888 335360 10940
rect 335412 10928 335418 10940
rect 392026 10928 392032 10940
rect 335412 10900 392032 10928
rect 335412 10888 335418 10900
rect 392026 10888 392032 10900
rect 392084 10888 392090 10940
rect 229370 10820 229376 10872
rect 229428 10860 229434 10872
rect 293954 10860 293960 10872
rect 229428 10832 293960 10860
rect 229428 10820 229434 10832
rect 293954 10820 293960 10832
rect 294012 10820 294018 10872
rect 381538 10820 381544 10872
rect 381596 10860 381602 10872
rect 442994 10860 443000 10872
rect 381596 10832 443000 10860
rect 381596 10820 381602 10832
rect 442994 10820 443000 10832
rect 443052 10820 443058 10872
rect 180242 10752 180248 10804
rect 180300 10792 180306 10804
rect 280246 10792 280252 10804
rect 180300 10764 280252 10792
rect 180300 10752 180306 10764
rect 280246 10752 280252 10764
rect 280304 10752 280310 10804
rect 338206 10752 338212 10804
rect 338264 10792 338270 10804
rect 403526 10792 403532 10804
rect 338264 10764 403532 10792
rect 338264 10752 338270 10764
rect 403526 10752 403532 10764
rect 403584 10752 403590 10804
rect 403710 10752 403716 10804
rect 403768 10792 403774 10804
rect 445754 10792 445760 10804
rect 403768 10764 445760 10792
rect 403768 10752 403774 10764
rect 445754 10752 445760 10764
rect 445812 10752 445818 10804
rect 172698 10684 172704 10736
rect 172756 10724 172762 10736
rect 278774 10724 278780 10736
rect 172756 10696 278780 10724
rect 172756 10684 172762 10696
rect 278774 10684 278780 10696
rect 278832 10684 278838 10736
rect 339586 10684 339592 10736
rect 339644 10724 339650 10736
rect 407206 10724 407212 10736
rect 339644 10696 407212 10724
rect 339644 10684 339650 10696
rect 407206 10684 407212 10696
rect 407264 10684 407270 10736
rect 168374 10616 168380 10668
rect 168432 10656 168438 10668
rect 277486 10656 277492 10668
rect 168432 10628 277492 10656
rect 168432 10616 168438 10628
rect 277486 10616 277492 10628
rect 277544 10616 277550 10668
rect 339494 10616 339500 10668
rect 339552 10656 339558 10668
rect 410794 10656 410800 10668
rect 339552 10628 410800 10656
rect 339552 10616 339558 10628
rect 410794 10616 410800 10628
rect 410852 10616 410858 10668
rect 166074 10548 166080 10600
rect 166132 10588 166138 10600
rect 277578 10588 277584 10600
rect 166132 10560 277584 10588
rect 166132 10548 166138 10560
rect 277578 10548 277584 10560
rect 277636 10548 277642 10600
rect 301498 10548 301504 10600
rect 301556 10588 301562 10600
rect 425698 10588 425704 10600
rect 301556 10560 425704 10588
rect 301556 10548 301562 10560
rect 425698 10548 425704 10560
rect 425756 10548 425762 10600
rect 269758 10480 269764 10532
rect 269816 10520 269822 10532
rect 411254 10520 411260 10532
rect 269816 10492 411260 10520
rect 269816 10480 269822 10492
rect 411254 10480 411260 10492
rect 411312 10480 411318 10532
rect 77386 10412 77392 10464
rect 77444 10452 77450 10464
rect 103514 10452 103520 10464
rect 77444 10424 103520 10452
rect 77444 10412 77450 10424
rect 103514 10412 103520 10424
rect 103572 10412 103578 10464
rect 162026 10412 162032 10464
rect 162084 10452 162090 10464
rect 276014 10452 276020 10464
rect 162084 10424 276020 10452
rect 162084 10412 162090 10424
rect 276014 10412 276020 10424
rect 276072 10412 276078 10464
rect 283098 10412 283104 10464
rect 283156 10452 283162 10464
rect 306558 10452 306564 10464
rect 283156 10424 306564 10452
rect 283156 10412 283162 10424
rect 306558 10412 306564 10424
rect 306616 10412 306622 10464
rect 371234 10412 371240 10464
rect 371292 10452 371298 10464
rect 531406 10452 531412 10464
rect 371292 10424 531412 10452
rect 371292 10412 371298 10424
rect 531406 10412 531412 10424
rect 531464 10412 531470 10464
rect 33594 10344 33600 10396
rect 33652 10384 33658 10396
rect 62114 10384 62120 10396
rect 33652 10356 62120 10384
rect 33652 10344 33658 10356
rect 62114 10344 62120 10356
rect 62172 10344 62178 10396
rect 78674 10344 78680 10396
rect 78732 10384 78738 10396
rect 97442 10384 97448 10396
rect 78732 10356 97448 10384
rect 78732 10344 78738 10356
rect 97442 10344 97448 10356
rect 97500 10344 97506 10396
rect 103330 10344 103336 10396
rect 103388 10384 103394 10396
rect 139486 10384 139492 10396
rect 103388 10356 139492 10384
rect 103388 10344 103394 10356
rect 139486 10344 139492 10356
rect 139544 10344 139550 10396
rect 238754 10344 238760 10396
rect 238812 10384 238818 10396
rect 469858 10384 469864 10396
rect 238812 10356 469864 10384
rect 238812 10344 238818 10356
rect 469858 10344 469864 10356
rect 469916 10344 469922 10396
rect 478874 10344 478880 10396
rect 478932 10384 478938 10396
rect 499574 10384 499580 10396
rect 478932 10356 499580 10384
rect 478932 10344 478938 10356
rect 499574 10344 499580 10356
rect 499632 10344 499638 10396
rect 56778 10276 56784 10328
rect 56836 10316 56842 10328
rect 126238 10316 126244 10328
rect 56836 10288 126244 10316
rect 56836 10276 56842 10288
rect 126238 10276 126244 10288
rect 126296 10276 126302 10328
rect 240134 10276 240140 10328
rect 240192 10316 240198 10328
rect 476482 10316 476488 10328
rect 240192 10288 476488 10316
rect 240192 10276 240198 10288
rect 476482 10276 476488 10288
rect 476540 10276 476546 10328
rect 483106 10276 483112 10328
rect 483164 10316 483170 10328
rect 517882 10316 517888 10328
rect 483164 10288 517888 10316
rect 483164 10276 483170 10288
rect 517882 10276 517888 10288
rect 517940 10276 517946 10328
rect 400674 9528 400680 9580
rect 400732 9568 400738 9580
rect 444374 9568 444380 9580
rect 400732 9540 444380 9568
rect 400732 9528 400738 9540
rect 444374 9528 444380 9540
rect 444432 9528 444438 9580
rect 254670 9460 254676 9512
rect 254728 9500 254734 9512
rect 298738 9500 298744 9512
rect 254728 9472 298744 9500
rect 254728 9460 254734 9472
rect 298738 9460 298744 9472
rect 298796 9460 298802 9512
rect 356698 9460 356704 9512
rect 356756 9500 356762 9512
rect 471054 9500 471060 9512
rect 356756 9472 471060 9500
rect 356756 9460 356762 9472
rect 471054 9460 471060 9472
rect 471112 9460 471118 9512
rect 291378 9392 291384 9444
rect 291436 9432 291442 9444
rect 421558 9432 421564 9444
rect 291436 9404 421564 9432
rect 291436 9392 291442 9404
rect 421558 9392 421564 9404
rect 421616 9392 421622 9444
rect 190822 9324 190828 9376
rect 190880 9364 190886 9376
rect 283006 9364 283012 9376
rect 190880 9336 283012 9364
rect 190880 9324 190886 9336
rect 283006 9324 283012 9336
rect 283064 9324 283070 9376
rect 368474 9324 368480 9376
rect 368532 9364 368538 9376
rect 524230 9364 524236 9376
rect 368532 9336 524236 9364
rect 368532 9324 368538 9336
rect 524230 9324 524236 9336
rect 524288 9324 524294 9376
rect 222286 9256 222292 9308
rect 222344 9296 222350 9308
rect 402514 9296 402520 9308
rect 222344 9268 402520 9296
rect 222344 9256 222350 9268
rect 402514 9256 402520 9268
rect 402572 9256 402578 9308
rect 222194 9188 222200 9240
rect 222252 9228 222258 9240
rect 406010 9228 406016 9240
rect 222252 9200 406016 9228
rect 222252 9188 222258 9200
rect 406010 9188 406016 9200
rect 406068 9188 406074 9240
rect 223574 9120 223580 9172
rect 223632 9160 223638 9172
rect 409598 9160 409604 9172
rect 223632 9132 409604 9160
rect 223632 9120 223638 9132
rect 409598 9120 409604 9132
rect 409656 9120 409662 9172
rect 79318 9052 79324 9104
rect 79376 9092 79382 9104
rect 90358 9092 90364 9104
rect 79376 9064 90364 9092
rect 79376 9052 79382 9064
rect 90358 9052 90364 9064
rect 90416 9052 90422 9104
rect 95142 9052 95148 9104
rect 95200 9092 95206 9104
rect 107746 9092 107752 9104
rect 95200 9064 107752 9092
rect 95200 9052 95206 9064
rect 107746 9052 107752 9064
rect 107804 9052 107810 9104
rect 226334 9052 226340 9104
rect 226392 9092 226398 9104
rect 420178 9092 420184 9104
rect 226392 9064 420184 9092
rect 226392 9052 226398 9064
rect 420178 9052 420184 9064
rect 420236 9052 420242 9104
rect 56042 8984 56048 9036
rect 56100 9024 56106 9036
rect 97994 9024 98000 9036
rect 56100 8996 98000 9024
rect 56100 8984 56106 8996
rect 97994 8984 98000 8996
rect 98052 8984 98058 9036
rect 164326 8984 164332 9036
rect 164384 9024 164390 9036
rect 179046 9024 179052 9036
rect 164384 8996 179052 9024
rect 164384 8984 164390 8996
rect 179046 8984 179052 8996
rect 179104 8984 179110 9036
rect 227806 8984 227812 9036
rect 227864 9024 227870 9036
rect 423766 9024 423772 9036
rect 227864 8996 423772 9024
rect 227864 8984 227870 8996
rect 423766 8984 423772 8996
rect 423824 8984 423830 9036
rect 424318 8984 424324 9036
rect 424376 9024 424382 9036
rect 480530 9024 480536 9036
rect 424376 8996 480536 9024
rect 424376 8984 424382 8996
rect 480530 8984 480536 8996
rect 480588 8984 480594 9036
rect 482278 8984 482284 9036
rect 482336 9024 482342 9036
rect 497090 9024 497096 9036
rect 482336 8996 497096 9024
rect 482336 8984 482342 8996
rect 497090 8984 497096 8996
rect 497148 8984 497154 9036
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 57974 8956 57980 8968
rect 12400 8928 57980 8956
rect 12400 8916 12406 8928
rect 57974 8916 57980 8928
rect 58032 8916 58038 8968
rect 71498 8916 71504 8968
rect 71556 8956 71562 8968
rect 130378 8956 130384 8968
rect 71556 8928 130384 8956
rect 71556 8916 71562 8928
rect 130378 8916 130384 8928
rect 130436 8916 130442 8968
rect 173158 8916 173164 8968
rect 173216 8956 173222 8968
rect 203886 8956 203892 8968
rect 173216 8928 203892 8956
rect 173216 8916 173222 8928
rect 203886 8916 203892 8928
rect 203944 8916 203950 8968
rect 230474 8916 230480 8968
rect 230532 8956 230538 8968
rect 437934 8956 437940 8968
rect 230532 8928 437940 8956
rect 230532 8916 230538 8928
rect 437934 8916 437940 8928
rect 437992 8916 437998 8968
rect 483014 8916 483020 8968
rect 483072 8956 483078 8968
rect 514754 8956 514760 8968
rect 483072 8928 514760 8956
rect 483072 8916 483078 8928
rect 514754 8916 514760 8928
rect 514812 8916 514818 8968
rect 428458 8304 428464 8356
rect 428516 8344 428522 8356
rect 434438 8344 434444 8356
rect 428516 8316 434444 8344
rect 428516 8304 428522 8316
rect 434438 8304 434444 8316
rect 434496 8304 434502 8356
rect 74626 8236 74632 8288
rect 74684 8276 74690 8288
rect 83274 8276 83280 8288
rect 74684 8248 83280 8276
rect 74684 8236 74690 8248
rect 83274 8236 83280 8248
rect 83332 8236 83338 8288
rect 224218 8236 224224 8288
rect 224276 8276 224282 8288
rect 225138 8276 225144 8288
rect 224276 8248 225144 8276
rect 224276 8236 224282 8248
rect 225138 8236 225144 8248
rect 225196 8236 225202 8288
rect 258258 8236 258264 8288
rect 258316 8276 258322 8288
rect 300118 8276 300124 8288
rect 258316 8248 300124 8276
rect 258316 8236 258322 8248
rect 300118 8236 300124 8248
rect 300176 8236 300182 8288
rect 332594 8236 332600 8288
rect 332652 8276 332658 8288
rect 382366 8276 382372 8288
rect 332652 8248 382372 8276
rect 332652 8236 332658 8248
rect 382366 8236 382372 8248
rect 382424 8236 382430 8288
rect 244090 8168 244096 8220
rect 244148 8208 244154 8220
rect 296806 8208 296812 8220
rect 244148 8180 296812 8208
rect 244148 8168 244154 8180
rect 296806 8168 296812 8180
rect 296864 8168 296870 8220
rect 333974 8168 333980 8220
rect 334032 8208 334038 8220
rect 385954 8208 385960 8220
rect 334032 8180 385960 8208
rect 334032 8168 334038 8180
rect 385954 8168 385960 8180
rect 386012 8168 386018 8220
rect 282086 8100 282092 8152
rect 282144 8140 282150 8152
rect 422294 8140 422300 8152
rect 282144 8112 422300 8140
rect 282144 8100 282150 8112
rect 422294 8100 422300 8112
rect 422352 8100 422358 8152
rect 242158 8032 242164 8084
rect 242216 8072 242222 8084
rect 303154 8072 303160 8084
rect 242216 8044 303160 8072
rect 242216 8032 242222 8044
rect 303154 8032 303160 8044
rect 303212 8032 303218 8084
rect 375374 8032 375380 8084
rect 375432 8072 375438 8084
rect 549070 8072 549076 8084
rect 375432 8044 549076 8072
rect 375432 8032 375438 8044
rect 549070 8032 549076 8044
rect 549128 8032 549134 8084
rect 199378 7964 199384 8016
rect 199436 8004 199442 8016
rect 274818 8004 274824 8016
rect 199436 7976 274824 8004
rect 199436 7964 199442 7976
rect 274818 7964 274824 7976
rect 274876 7964 274882 8016
rect 376846 7964 376852 8016
rect 376904 8004 376910 8016
rect 552658 8004 552664 8016
rect 376904 7976 552664 8004
rect 376904 7964 376910 7976
rect 552658 7964 552664 7976
rect 552716 7964 552722 8016
rect 205082 7896 205088 7948
rect 205140 7936 205146 7948
rect 287054 7936 287060 7948
rect 205140 7908 287060 7936
rect 205140 7896 205146 7908
rect 287054 7896 287060 7908
rect 287112 7896 287118 7948
rect 328546 7896 328552 7948
rect 328604 7936 328610 7948
rect 368198 7936 368204 7948
rect 328604 7908 368204 7936
rect 328604 7896 328610 7908
rect 368198 7896 368204 7908
rect 368256 7896 368262 7948
rect 376938 7896 376944 7948
rect 376996 7936 377002 7948
rect 556154 7936 556160 7948
rect 376996 7908 556160 7936
rect 376996 7896 377002 7908
rect 556154 7896 556160 7908
rect 556212 7896 556218 7948
rect 187326 7828 187332 7880
rect 187384 7868 187390 7880
rect 282178 7868 282184 7880
rect 187384 7840 282184 7868
rect 187384 7828 187390 7840
rect 282178 7828 282184 7840
rect 282236 7828 282242 7880
rect 329834 7828 329840 7880
rect 329892 7868 329898 7880
rect 371694 7868 371700 7880
rect 329892 7840 371700 7868
rect 329892 7828 329898 7840
rect 371694 7828 371700 7840
rect 371752 7828 371758 7880
rect 378134 7828 378140 7880
rect 378192 7868 378198 7880
rect 559742 7868 559748 7880
rect 378192 7840 559748 7868
rect 378192 7828 378198 7840
rect 559742 7828 559748 7840
rect 559800 7828 559806 7880
rect 176746 7760 176752 7812
rect 176804 7800 176810 7812
rect 280154 7800 280160 7812
rect 176804 7772 280160 7800
rect 176804 7760 176810 7772
rect 280154 7760 280160 7772
rect 280212 7760 280218 7812
rect 297266 7760 297272 7812
rect 297324 7800 297330 7812
rect 310514 7800 310520 7812
rect 297324 7772 310520 7800
rect 297324 7760 297330 7772
rect 310514 7760 310520 7772
rect 310572 7760 310578 7812
rect 331214 7760 331220 7812
rect 331272 7800 331278 7812
rect 375282 7800 375288 7812
rect 331272 7772 375288 7800
rect 331272 7760 331278 7772
rect 375282 7760 375288 7772
rect 375340 7760 375346 7812
rect 380894 7760 380900 7812
rect 380952 7800 380958 7812
rect 570322 7800 570328 7812
rect 380952 7772 570328 7800
rect 380952 7760 380958 7772
rect 570322 7760 570328 7772
rect 570380 7760 570386 7812
rect 80054 7692 80060 7744
rect 80112 7732 80118 7744
rect 104526 7732 104532 7744
rect 80112 7704 104532 7732
rect 80112 7692 80118 7704
rect 104526 7692 104532 7704
rect 104584 7692 104590 7744
rect 200114 7692 200120 7744
rect 200172 7732 200178 7744
rect 320910 7732 320916 7744
rect 200172 7704 320916 7732
rect 200172 7692 200178 7704
rect 320910 7692 320916 7704
rect 320968 7692 320974 7744
rect 331306 7692 331312 7744
rect 331364 7732 331370 7744
rect 378870 7732 378876 7744
rect 331364 7704 378876 7732
rect 331364 7692 331370 7704
rect 378870 7692 378876 7704
rect 378928 7692 378934 7744
rect 382458 7692 382464 7744
rect 382516 7732 382522 7744
rect 573910 7732 573916 7744
rect 382516 7704 573916 7732
rect 382516 7692 382522 7704
rect 573910 7692 573916 7704
rect 573968 7692 573974 7744
rect 26510 7624 26516 7676
rect 26568 7664 26574 7676
rect 60734 7664 60740 7676
rect 26568 7636 60740 7664
rect 26568 7624 26574 7636
rect 60734 7624 60740 7636
rect 60792 7624 60798 7676
rect 62022 7624 62028 7676
rect 62080 7664 62086 7676
rect 70486 7664 70492 7676
rect 62080 7636 70492 7664
rect 62080 7624 62086 7636
rect 70486 7624 70492 7636
rect 70544 7624 70550 7676
rect 78582 7624 78588 7676
rect 78640 7664 78646 7676
rect 132494 7664 132500 7676
rect 78640 7636 132500 7664
rect 78640 7624 78646 7636
rect 132494 7624 132500 7636
rect 132552 7624 132558 7676
rect 136450 7624 136456 7676
rect 136508 7664 136514 7676
rect 153194 7664 153200 7676
rect 136508 7636 153200 7664
rect 136508 7624 136514 7636
rect 153194 7624 153200 7636
rect 153252 7624 153258 7676
rect 162946 7624 162952 7676
rect 163004 7664 163010 7676
rect 175458 7664 175464 7676
rect 163004 7636 175464 7664
rect 163004 7624 163010 7636
rect 175458 7624 175464 7636
rect 175516 7624 175522 7676
rect 175918 7624 175924 7676
rect 175976 7664 175982 7676
rect 189718 7664 189724 7676
rect 175976 7636 189724 7664
rect 175976 7624 175982 7636
rect 189718 7624 189724 7636
rect 189776 7624 189782 7676
rect 191098 7624 191104 7676
rect 191156 7664 191162 7676
rect 207382 7664 207388 7676
rect 191156 7636 207388 7664
rect 191156 7624 191162 7636
rect 207382 7624 207388 7636
rect 207440 7624 207446 7676
rect 209774 7624 209780 7676
rect 209832 7664 209838 7676
rect 356330 7664 356336 7676
rect 209832 7636 356336 7664
rect 209832 7624 209838 7636
rect 356330 7624 356336 7636
rect 356388 7624 356394 7676
rect 382274 7624 382280 7676
rect 382332 7664 382338 7676
rect 577406 7664 577412 7676
rect 382332 7636 577412 7664
rect 382332 7624 382338 7636
rect 577406 7624 577412 7636
rect 577464 7624 577470 7676
rect 38378 7556 38384 7608
rect 38436 7596 38442 7608
rect 93118 7596 93124 7608
rect 38436 7568 93124 7596
rect 38436 7556 38442 7568
rect 93118 7556 93124 7568
rect 93176 7556 93182 7608
rect 114646 7556 114652 7608
rect 114704 7596 114710 7608
rect 123478 7596 123484 7608
rect 114704 7568 123484 7596
rect 114704 7556 114710 7568
rect 123478 7556 123484 7568
rect 123536 7556 123542 7608
rect 131758 7556 131764 7608
rect 131816 7596 131822 7608
rect 385034 7596 385040 7608
rect 131816 7568 385040 7596
rect 131816 7556 131822 7568
rect 385034 7556 385040 7568
rect 385092 7556 385098 7608
rect 356054 7488 356060 7540
rect 356112 7528 356118 7540
rect 387794 7528 387800 7540
rect 356112 7500 387800 7528
rect 356112 7488 356118 7500
rect 387794 7488 387800 7500
rect 387852 7488 387858 7540
rect 279510 6808 279516 6860
rect 279568 6848 279574 6860
rect 306374 6848 306380 6860
rect 279568 6820 306380 6848
rect 279568 6808 279574 6820
rect 306374 6808 306380 6820
rect 306432 6808 306438 6860
rect 318794 6808 318800 6860
rect 318852 6848 318858 6860
rect 329190 6848 329196 6860
rect 318852 6820 329196 6848
rect 318852 6808 318858 6820
rect 329190 6808 329196 6820
rect 329248 6808 329254 6860
rect 337470 6808 337476 6860
rect 337528 6848 337534 6860
rect 403618 6848 403624 6860
rect 337528 6820 403624 6848
rect 337528 6808 337534 6820
rect 403618 6808 403624 6820
rect 403676 6808 403682 6860
rect 305178 6740 305184 6792
rect 305236 6780 305242 6792
rect 386414 6780 386420 6792
rect 305236 6752 386420 6780
rect 305236 6740 305242 6752
rect 386414 6740 386420 6752
rect 386472 6740 386478 6792
rect 266538 6672 266544 6724
rect 266596 6712 266602 6724
rect 367738 6712 367744 6724
rect 266596 6684 367744 6712
rect 266596 6672 266602 6684
rect 367738 6672 367744 6684
rect 367796 6672 367802 6724
rect 187694 6604 187700 6656
rect 187752 6644 187758 6656
rect 267734 6644 267740 6656
rect 187752 6616 267740 6644
rect 187752 6604 187758 6616
rect 267734 6604 267740 6616
rect 267792 6604 267798 6656
rect 276014 6604 276020 6656
rect 276072 6644 276078 6656
rect 305086 6644 305092 6656
rect 276072 6616 305092 6644
rect 276072 6604 276078 6616
rect 305086 6604 305092 6616
rect 305144 6604 305150 6656
rect 320174 6604 320180 6656
rect 320232 6644 320238 6656
rect 332686 6644 332692 6656
rect 320232 6616 332692 6644
rect 320232 6604 320238 6616
rect 332686 6604 332692 6616
rect 332744 6604 332750 6656
rect 357434 6604 357440 6656
rect 357492 6644 357498 6656
rect 481726 6644 481732 6656
rect 357492 6616 481732 6644
rect 357492 6604 357498 6616
rect 481726 6604 481732 6616
rect 481784 6604 481790 6656
rect 187786 6536 187792 6588
rect 187844 6576 187850 6588
rect 271230 6576 271236 6588
rect 187844 6548 271236 6576
rect 187844 6536 187850 6548
rect 271230 6536 271236 6548
rect 271288 6536 271294 6588
rect 272426 6536 272432 6588
rect 272484 6576 272490 6588
rect 304994 6576 305000 6588
rect 272484 6548 305000 6576
rect 272484 6536 272490 6548
rect 304994 6536 305000 6548
rect 305052 6536 305058 6588
rect 320266 6536 320272 6588
rect 320324 6576 320330 6588
rect 336274 6576 336280 6588
rect 320324 6548 336280 6576
rect 320324 6536 320330 6548
rect 336274 6536 336280 6548
rect 336332 6536 336338 6588
rect 358814 6536 358820 6588
rect 358872 6576 358878 6588
rect 485222 6576 485228 6588
rect 358872 6548 485228 6576
rect 358872 6536 358878 6548
rect 485222 6536 485228 6548
rect 485280 6536 485286 6588
rect 190454 6468 190460 6520
rect 190512 6508 190518 6520
rect 281902 6508 281908 6520
rect 190512 6480 281908 6508
rect 190512 6468 190518 6480
rect 281902 6468 281908 6480
rect 281960 6468 281966 6520
rect 321554 6468 321560 6520
rect 321612 6508 321618 6520
rect 339862 6508 339868 6520
rect 321612 6480 339868 6508
rect 321612 6468 321618 6480
rect 339862 6468 339868 6480
rect 339920 6468 339926 6520
rect 360194 6468 360200 6520
rect 360252 6508 360258 6520
rect 488810 6508 488816 6520
rect 360252 6480 488816 6508
rect 360252 6468 360258 6480
rect 488810 6468 488816 6480
rect 488868 6468 488874 6520
rect 191834 6400 191840 6452
rect 191892 6440 191898 6452
rect 285398 6440 285404 6452
rect 191892 6412 285404 6440
rect 191892 6400 191898 6412
rect 285398 6400 285404 6412
rect 285456 6400 285462 6452
rect 286594 6400 286600 6452
rect 286652 6440 286658 6452
rect 307754 6440 307760 6452
rect 286652 6412 307760 6440
rect 286652 6400 286658 6412
rect 307754 6400 307760 6412
rect 307812 6400 307818 6452
rect 322934 6400 322940 6452
rect 322992 6440 322998 6452
rect 343358 6440 343364 6452
rect 322992 6412 343364 6440
rect 322992 6400 322998 6412
rect 343358 6400 343364 6412
rect 343416 6400 343422 6452
rect 363046 6400 363052 6452
rect 363104 6440 363110 6452
rect 499390 6440 499396 6452
rect 363104 6412 499396 6440
rect 363104 6400 363110 6412
rect 499390 6400 499396 6412
rect 499448 6400 499454 6452
rect 191926 6332 191932 6384
rect 191984 6372 191990 6384
rect 288986 6372 288992 6384
rect 191984 6344 288992 6372
rect 191984 6332 191990 6344
rect 288986 6332 288992 6344
rect 289044 6332 289050 6384
rect 290182 6332 290188 6384
rect 290240 6372 290246 6384
rect 309134 6372 309140 6384
rect 290240 6344 309140 6372
rect 290240 6332 290246 6344
rect 309134 6332 309140 6344
rect 309192 6332 309198 6384
rect 323026 6332 323032 6384
rect 323084 6372 323090 6384
rect 346946 6372 346952 6384
rect 323084 6344 346952 6372
rect 323084 6332 323090 6344
rect 346946 6332 346952 6344
rect 347004 6332 347010 6384
rect 362954 6332 362960 6384
rect 363012 6372 363018 6384
rect 502978 6372 502984 6384
rect 363012 6344 502984 6372
rect 363012 6332 363018 6344
rect 502978 6332 502984 6344
rect 503036 6332 503042 6384
rect 91554 6264 91560 6316
rect 91612 6304 91618 6316
rect 106918 6304 106924 6316
rect 91612 6276 106924 6304
rect 91612 6264 91618 6276
rect 106918 6264 106924 6276
rect 106976 6264 106982 6316
rect 193214 6264 193220 6316
rect 193272 6304 193278 6316
rect 292574 6304 292580 6316
rect 193272 6276 292580 6304
rect 193272 6264 193278 6276
rect 292574 6264 292580 6276
rect 292632 6264 292638 6316
rect 293678 6264 293684 6316
rect 293736 6304 293742 6316
rect 309226 6304 309232 6316
rect 293736 6276 309232 6304
rect 293736 6264 293742 6276
rect 309226 6264 309232 6276
rect 309284 6264 309290 6316
rect 324314 6264 324320 6316
rect 324372 6304 324378 6316
rect 350442 6304 350448 6316
rect 324372 6276 350448 6304
rect 324372 6264 324378 6276
rect 350442 6264 350448 6276
rect 350500 6264 350506 6316
rect 364334 6264 364340 6316
rect 364392 6304 364398 6316
rect 506474 6304 506480 6316
rect 364392 6276 506480 6304
rect 364392 6264 364398 6276
rect 506474 6264 506480 6276
rect 506532 6264 506538 6316
rect 81434 6196 81440 6248
rect 81492 6236 81498 6248
rect 108114 6236 108120 6248
rect 81492 6208 108120 6236
rect 81492 6196 81498 6208
rect 108114 6196 108120 6208
rect 108172 6196 108178 6248
rect 129366 6196 129372 6248
rect 129424 6236 129430 6248
rect 151906 6236 151912 6248
rect 129424 6208 151912 6236
rect 129424 6196 129430 6208
rect 151906 6196 151912 6208
rect 151964 6196 151970 6248
rect 194686 6196 194692 6248
rect 194744 6236 194750 6248
rect 296070 6236 296076 6248
rect 194744 6208 296076 6236
rect 194744 6196 194750 6208
rect 296070 6196 296076 6208
rect 296128 6196 296134 6248
rect 327074 6196 327080 6248
rect 327132 6236 327138 6248
rect 361114 6236 361120 6248
rect 327132 6208 361120 6236
rect 327132 6196 327138 6208
rect 361114 6196 361120 6208
rect 361172 6196 361178 6248
rect 365714 6196 365720 6248
rect 365772 6236 365778 6248
rect 510062 6236 510068 6248
rect 365772 6208 510068 6236
rect 365772 6196 365778 6208
rect 510062 6196 510068 6208
rect 510120 6196 510126 6248
rect 512638 6196 512644 6248
rect 512696 6236 512702 6248
rect 525426 6236 525432 6248
rect 512696 6208 525432 6236
rect 512696 6196 512702 6208
rect 525426 6196 525432 6208
rect 525484 6196 525490 6248
rect 566 6128 572 6180
rect 624 6168 630 6180
rect 54478 6168 54484 6180
rect 624 6140 54484 6168
rect 624 6128 630 6140
rect 54478 6128 54484 6140
rect 54536 6128 54542 6180
rect 58434 6128 58440 6180
rect 58492 6168 58498 6180
rect 69198 6168 69204 6180
rect 58492 6140 69204 6168
rect 58492 6128 58498 6140
rect 69198 6128 69204 6140
rect 69256 6128 69262 6180
rect 76006 6128 76012 6180
rect 76064 6168 76070 6180
rect 86862 6168 86868 6180
rect 76064 6140 86868 6168
rect 76064 6128 76070 6140
rect 86862 6128 86868 6140
rect 86920 6128 86926 6180
rect 96246 6128 96252 6180
rect 96304 6168 96310 6180
rect 136634 6168 136640 6180
rect 96304 6140 136640 6168
rect 96304 6128 96310 6140
rect 136634 6128 136640 6140
rect 136692 6128 136698 6180
rect 165614 6128 165620 6180
rect 165672 6168 165678 6180
rect 182542 6168 182548 6180
rect 165672 6140 182548 6168
rect 165672 6128 165678 6140
rect 182542 6128 182548 6140
rect 182600 6128 182606 6180
rect 194778 6128 194784 6180
rect 194836 6168 194842 6180
rect 299658 6168 299664 6180
rect 194836 6140 299664 6168
rect 194836 6128 194842 6140
rect 299658 6128 299664 6140
rect 299716 6128 299722 6180
rect 304350 6128 304356 6180
rect 304408 6168 304414 6180
rect 311894 6168 311900 6180
rect 304408 6140 311900 6168
rect 304408 6128 304414 6140
rect 311894 6128 311900 6140
rect 311952 6128 311958 6180
rect 328454 6128 328460 6180
rect 328512 6168 328518 6180
rect 364610 6168 364616 6180
rect 328512 6140 364616 6168
rect 328512 6128 328518 6140
rect 364610 6128 364616 6140
rect 364668 6128 364674 6180
rect 365806 6128 365812 6180
rect 365864 6168 365870 6180
rect 513558 6168 513564 6180
rect 365864 6140 513564 6168
rect 365864 6128 365870 6140
rect 513558 6128 513564 6140
rect 513616 6128 513622 6180
rect 317414 5584 317420 5636
rect 317472 5624 317478 5636
rect 325602 5624 325608 5636
rect 317472 5596 325608 5624
rect 317472 5584 317478 5596
rect 325602 5584 325608 5596
rect 325660 5584 325666 5636
rect 74534 5516 74540 5568
rect 74592 5556 74598 5568
rect 79686 5556 79692 5568
rect 74592 5528 79692 5556
rect 74592 5516 74598 5528
rect 79686 5516 79692 5528
rect 79744 5516 79750 5568
rect 114554 5516 114560 5568
rect 114612 5556 114618 5568
rect 119890 5556 119896 5568
rect 114612 5528 119896 5556
rect 114612 5516 114618 5528
rect 119890 5516 119896 5528
rect 119948 5516 119954 5568
rect 184198 5516 184204 5568
rect 184256 5556 184262 5568
rect 186130 5556 186136 5568
rect 184256 5528 186136 5556
rect 184256 5516 184262 5528
rect 186130 5516 186136 5528
rect 186188 5516 186194 5568
rect 307938 5516 307944 5568
rect 307996 5556 308002 5568
rect 313366 5556 313372 5568
rect 307996 5528 313372 5556
rect 307996 5516 308002 5528
rect 313366 5516 313372 5528
rect 313424 5516 313430 5568
rect 317506 5516 317512 5568
rect 317564 5556 317570 5568
rect 322106 5556 322112 5568
rect 317564 5528 322112 5556
rect 317564 5516 317570 5528
rect 322106 5516 322112 5528
rect 322164 5516 322170 5568
rect 246298 5380 246304 5432
rect 246356 5420 246362 5432
rect 257062 5420 257068 5432
rect 246356 5392 257068 5420
rect 246356 5380 246362 5392
rect 257062 5380 257068 5392
rect 257120 5380 257126 5432
rect 178034 5312 178040 5364
rect 178092 5352 178098 5364
rect 232222 5352 232228 5364
rect 178092 5324 232228 5352
rect 178092 5312 178098 5324
rect 232222 5312 232228 5324
rect 232280 5312 232286 5364
rect 240502 5312 240508 5364
rect 240560 5352 240566 5364
rect 295978 5352 295984 5364
rect 240560 5324 295984 5352
rect 240560 5312 240566 5324
rect 295978 5312 295984 5324
rect 296036 5312 296042 5364
rect 348050 5312 348056 5364
rect 348108 5352 348114 5364
rect 418798 5352 418804 5364
rect 348108 5324 418804 5352
rect 348108 5312 348114 5324
rect 418798 5312 418804 5324
rect 418856 5312 418862 5364
rect 201586 5244 201592 5296
rect 201644 5284 201650 5296
rect 285674 5284 285680 5296
rect 201644 5256 285680 5284
rect 201644 5244 201650 5256
rect 285674 5244 285680 5256
rect 285732 5244 285738 5296
rect 317322 5244 317328 5296
rect 317380 5284 317386 5296
rect 429286 5284 429292 5296
rect 317380 5256 429292 5284
rect 317380 5244 317386 5256
rect 429286 5244 429292 5256
rect 429344 5244 429350 5296
rect 54938 5176 54944 5228
rect 54996 5216 55002 5228
rect 67634 5216 67640 5228
rect 54996 5188 67640 5216
rect 54996 5176 55002 5188
rect 67634 5176 67640 5188
rect 67692 5176 67698 5228
rect 223942 5176 223948 5228
rect 224000 5216 224006 5228
rect 407758 5216 407764 5228
rect 224000 5188 407764 5216
rect 224000 5176 224006 5188
rect 407758 5176 407764 5188
rect 407816 5176 407822 5228
rect 52546 5108 52552 5160
rect 52604 5148 52610 5160
rect 96706 5148 96712 5160
rect 52604 5120 96712 5148
rect 52604 5108 52610 5120
rect 96706 5108 96712 5120
rect 96764 5108 96770 5160
rect 231854 5108 231860 5160
rect 231912 5148 231918 5160
rect 445018 5148 445024 5160
rect 231912 5120 445024 5148
rect 231912 5108 231918 5120
rect 445018 5108 445024 5120
rect 445076 5108 445082 5160
rect 48958 5040 48964 5092
rect 49016 5080 49022 5092
rect 96614 5080 96620 5092
rect 49016 5052 96620 5080
rect 49016 5040 49022 5052
rect 96614 5040 96620 5052
rect 96672 5040 96678 5092
rect 175274 5040 175280 5092
rect 175332 5080 175338 5092
rect 221550 5080 221556 5092
rect 175332 5052 221556 5080
rect 175332 5040 175338 5052
rect 221550 5040 221556 5052
rect 221608 5040 221614 5092
rect 249794 5040 249800 5092
rect 249852 5080 249858 5092
rect 512454 5080 512460 5092
rect 249852 5052 512460 5080
rect 249852 5040 249858 5052
rect 512454 5040 512460 5052
rect 512512 5040 512518 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 56594 5012 56600 5024
rect 7708 4984 56600 5012
rect 7708 4972 7714 4984
rect 56594 4972 56600 4984
rect 56652 4972 56658 5024
rect 82814 4972 82820 5024
rect 82872 5012 82878 5024
rect 115198 5012 115204 5024
rect 82872 4984 115204 5012
rect 82872 4972 82878 4984
rect 115198 4972 115204 4984
rect 115256 4972 115262 5024
rect 179414 4972 179420 5024
rect 179472 5012 179478 5024
rect 235810 5012 235816 5024
rect 179472 4984 235816 5012
rect 179472 4972 179478 4984
rect 235810 4972 235816 4984
rect 235868 4972 235874 5024
rect 255314 4972 255320 5024
rect 255372 5012 255378 5024
rect 533706 5012 533712 5024
rect 255372 4984 533712 5012
rect 255372 4972 255378 4984
rect 533706 4972 533712 4984
rect 533764 4972 533770 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 56686 4944 56692 4956
rect 2924 4916 56692 4944
rect 2924 4904 2930 4916
rect 56686 4904 56692 4916
rect 56744 4904 56750 4956
rect 85850 4904 85856 4956
rect 85908 4944 85914 4956
rect 122282 4944 122288 4956
rect 85908 4916 122288 4944
rect 85908 4904 85914 4916
rect 122282 4904 122288 4916
rect 122340 4904 122346 4956
rect 179506 4904 179512 4956
rect 179564 4944 179570 4956
rect 239306 4944 239312 4956
rect 179564 4916 239312 4944
rect 179564 4904 179570 4916
rect 239306 4904 239312 4916
rect 239364 4904 239370 4956
rect 256694 4904 256700 4956
rect 256752 4944 256758 4956
rect 537202 4944 537208 4956
rect 256752 4916 537208 4944
rect 256752 4904 256758 4916
rect 537202 4904 537208 4916
rect 537260 4904 537266 4956
rect 8754 4836 8760 4888
rect 8812 4876 8818 4888
rect 86954 4876 86960 4888
rect 8812 4848 86960 4876
rect 8812 4836 8818 4848
rect 86954 4836 86960 4848
rect 87012 4836 87018 4888
rect 170398 4836 170404 4888
rect 170456 4876 170462 4888
rect 171962 4876 171968 4888
rect 170456 4848 171968 4876
rect 170456 4836 170462 4848
rect 171962 4836 171968 4848
rect 172020 4836 172026 4888
rect 182266 4836 182272 4888
rect 182324 4876 182330 4888
rect 246390 4876 246396 4888
rect 182324 4848 246396 4876
rect 182324 4836 182330 4848
rect 246390 4836 246396 4848
rect 246448 4836 246454 4888
rect 256786 4836 256792 4888
rect 256844 4876 256850 4888
rect 540790 4876 540796 4888
rect 256844 4848 540796 4876
rect 256844 4836 256850 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 85666 4808 85672 4820
rect 4120 4780 85672 4808
rect 4120 4768 4126 4780
rect 85666 4768 85672 4780
rect 85724 4768 85730 4820
rect 125870 4768 125876 4820
rect 125928 4808 125934 4820
rect 150710 4808 150716 4820
rect 125928 4780 150716 4808
rect 125928 4768 125934 4780
rect 150710 4768 150716 4780
rect 150768 4768 150774 4820
rect 182174 4768 182180 4820
rect 182232 4808 182238 4820
rect 249978 4808 249984 4820
rect 182232 4780 249984 4808
rect 182232 4768 182238 4780
rect 249978 4768 249984 4780
rect 250036 4768 250042 4820
rect 258074 4768 258080 4820
rect 258132 4808 258138 4820
rect 544378 4808 544384 4820
rect 258132 4780 544384 4808
rect 258132 4768 258138 4780
rect 544378 4768 544384 4780
rect 544436 4768 544442 4820
rect 569218 4768 569224 4820
rect 569276 4808 569282 4820
rect 579798 4808 579804 4820
rect 569276 4780 579804 4808
rect 569276 4768 569282 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 65518 4156 65524 4208
rect 65576 4196 65582 4208
rect 70394 4196 70400 4208
rect 65576 4168 70400 4196
rect 65576 4156 65582 4168
rect 70394 4156 70400 4168
rect 70452 4156 70458 4208
rect 161474 4156 161480 4208
rect 161532 4196 161538 4208
rect 168466 4196 168472 4208
rect 161532 4168 168472 4196
rect 161532 4156 161538 4168
rect 168466 4156 168472 4168
rect 168524 4156 168530 4208
rect 448606 4156 448612 4208
rect 448664 4196 448670 4208
rect 449986 4196 449992 4208
rect 448664 4168 449992 4196
rect 448664 4156 448670 4168
rect 449986 4156 449992 4168
rect 450044 4156 450050 4208
rect 46658 4088 46664 4140
rect 46716 4128 46722 4140
rect 124214 4128 124220 4140
rect 46716 4100 124220 4128
rect 46716 4088 46722 4100
rect 124214 4088 124220 4100
rect 124272 4088 124278 4140
rect 376478 4088 376484 4140
rect 376536 4128 376542 4140
rect 385678 4128 385684 4140
rect 376536 4100 385684 4128
rect 376536 4088 376542 4100
rect 385678 4088 385684 4100
rect 385736 4088 385742 4140
rect 422570 4088 422576 4140
rect 422628 4128 422634 4140
rect 459646 4128 459652 4140
rect 422628 4100 459652 4128
rect 422628 4088 422634 4100
rect 459646 4088 459652 4100
rect 459704 4088 459710 4140
rect 491294 4088 491300 4140
rect 491352 4128 491358 4140
rect 550266 4128 550272 4140
rect 491352 4100 550272 4128
rect 491352 4088 491358 4100
rect 550266 4088 550272 4100
rect 550324 4088 550330 4140
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 122926 4060 122932 4072
rect 43128 4032 122932 4060
rect 43128 4020 43134 4032
rect 122926 4020 122932 4032
rect 122984 4020 122990 4072
rect 362310 4020 362316 4072
rect 362368 4060 362374 4072
rect 378778 4060 378784 4072
rect 362368 4032 378784 4060
rect 362368 4020 362374 4032
rect 378778 4020 378784 4032
rect 378836 4020 378842 4072
rect 411898 4060 411904 4072
rect 393286 4032 411904 4060
rect 39574 3952 39580 4004
rect 39632 3992 39638 4004
rect 122834 3992 122840 4004
rect 39632 3964 122840 3992
rect 39632 3952 39638 3964
rect 122834 3952 122840 3964
rect 122892 3952 122898 4004
rect 333882 3952 333888 4004
rect 333940 3992 333946 4004
rect 342898 3992 342904 4004
rect 333940 3964 342904 3992
rect 333940 3952 333946 3964
rect 342898 3952 342904 3964
rect 342956 3952 342962 4004
rect 355226 3952 355232 4004
rect 355284 3992 355290 4004
rect 376018 3992 376024 4004
rect 355284 3964 376024 3992
rect 355284 3952 355290 3964
rect 376018 3952 376024 3964
rect 376076 3952 376082 4004
rect 379974 3952 379980 4004
rect 380032 3992 380038 4004
rect 393286 3992 393314 4032
rect 411898 4020 411904 4032
rect 411956 4020 411962 4072
rect 418982 4020 418988 4072
rect 419040 4060 419046 4072
rect 458174 4060 458180 4072
rect 419040 4032 458180 4060
rect 419040 4020 419046 4032
rect 458174 4020 458180 4032
rect 458232 4020 458238 4072
rect 492766 4020 492772 4072
rect 492824 4060 492830 4072
rect 553762 4060 553768 4072
rect 492824 4032 553768 4060
rect 492824 4020 492830 4032
rect 553762 4020 553768 4032
rect 553820 4020 553826 4072
rect 380032 3964 393314 3992
rect 380032 3952 380038 3964
rect 415486 3952 415492 4004
rect 415544 3992 415550 4004
rect 456794 3992 456800 4004
rect 415544 3964 456800 3992
rect 415544 3952 415550 3964
rect 456794 3952 456800 3964
rect 456852 3952 456858 4004
rect 494146 3952 494152 4004
rect 494204 3992 494210 4004
rect 557350 3992 557356 4004
rect 494204 3964 557356 3992
rect 494204 3952 494210 3964
rect 557350 3952 557356 3964
rect 557408 3952 557414 4004
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 121546 3924 121552 3936
rect 36044 3896 121552 3924
rect 36044 3884 36050 3896
rect 121546 3884 121552 3896
rect 121604 3884 121610 3936
rect 140038 3884 140044 3936
rect 140096 3924 140102 3936
rect 154758 3924 154764 3936
rect 140096 3896 154764 3924
rect 140096 3884 140102 3896
rect 154758 3884 154764 3896
rect 154816 3884 154822 3936
rect 251174 3884 251180 3936
rect 251232 3924 251238 3936
rect 252370 3924 252376 3936
rect 251232 3896 252376 3924
rect 251232 3884 251238 3896
rect 252370 3884 252376 3896
rect 252428 3884 252434 3936
rect 262950 3884 262956 3936
rect 263008 3924 263014 3936
rect 273898 3924 273904 3936
rect 263008 3896 273904 3924
rect 263008 3884 263014 3896
rect 273898 3884 273904 3896
rect 273956 3884 273962 3936
rect 305546 3884 305552 3936
rect 305604 3924 305610 3936
rect 312538 3924 312544 3936
rect 305604 3896 312544 3924
rect 305604 3884 305610 3896
rect 312538 3884 312544 3896
rect 312596 3884 312602 3936
rect 319714 3884 319720 3936
rect 319772 3924 319778 3936
rect 330478 3924 330484 3936
rect 319772 3896 330484 3924
rect 319772 3884 319778 3896
rect 330478 3884 330484 3896
rect 330536 3884 330542 3936
rect 340966 3884 340972 3936
rect 341024 3924 341030 3936
rect 353938 3924 353944 3936
rect 341024 3896 353944 3924
rect 341024 3884 341030 3896
rect 353938 3884 353944 3896
rect 353996 3884 354002 3936
rect 372890 3884 372896 3936
rect 372948 3924 372954 3936
rect 404998 3924 405004 3936
rect 372948 3896 405004 3924
rect 372948 3884 372954 3896
rect 404998 3884 405004 3896
rect 405056 3884 405062 3936
rect 411898 3884 411904 3936
rect 411956 3924 411962 3936
rect 456978 3924 456984 3936
rect 411956 3896 456984 3924
rect 411956 3884 411962 3896
rect 456978 3884 456984 3896
rect 457036 3884 457042 3936
rect 494054 3884 494060 3936
rect 494112 3924 494118 3936
rect 560846 3924 560852 3936
rect 494112 3896 560852 3924
rect 494112 3884 494118 3896
rect 560846 3884 560852 3896
rect 560904 3884 560910 3936
rect 32398 3816 32404 3868
rect 32456 3856 32462 3868
rect 120166 3856 120172 3868
rect 32456 3828 120172 3856
rect 32456 3816 32462 3828
rect 120166 3816 120172 3828
rect 120224 3816 120230 3868
rect 124674 3816 124680 3868
rect 124732 3856 124738 3868
rect 145006 3856 145012 3868
rect 124732 3828 145012 3856
rect 124732 3816 124738 3828
rect 145006 3816 145012 3828
rect 145064 3816 145070 3868
rect 176654 3816 176660 3868
rect 176712 3856 176718 3868
rect 177850 3856 177856 3868
rect 176712 3828 177856 3856
rect 176712 3816 176718 3828
rect 177850 3816 177856 3828
rect 177908 3816 177914 3868
rect 193214 3816 193220 3868
rect 193272 3856 193278 3868
rect 193398 3856 193404 3868
rect 193272 3828 193404 3856
rect 193272 3816 193278 3828
rect 193398 3816 193404 3828
rect 193456 3816 193462 3868
rect 209866 3816 209872 3868
rect 209924 3856 209930 3868
rect 210970 3856 210976 3868
rect 209924 3828 210976 3856
rect 209924 3816 209930 3828
rect 210970 3816 210976 3828
rect 211028 3816 211034 3868
rect 226426 3816 226432 3868
rect 226484 3856 226490 3868
rect 227530 3856 227536 3868
rect 226484 3828 227536 3856
rect 226484 3816 226490 3828
rect 227530 3816 227536 3828
rect 227588 3816 227594 3868
rect 234614 3816 234620 3868
rect 234672 3856 234678 3868
rect 269758 3856 269764 3868
rect 234672 3828 269764 3856
rect 234672 3816 234678 3828
rect 269758 3816 269764 3828
rect 269816 3816 269822 3868
rect 277118 3816 277124 3868
rect 277176 3856 277182 3868
rect 282086 3856 282092 3868
rect 277176 3828 282092 3856
rect 277176 3816 277182 3828
rect 282086 3816 282092 3828
rect 282144 3816 282150 3868
rect 287790 3816 287796 3868
rect 287848 3856 287854 3868
rect 294598 3856 294604 3868
rect 287848 3828 294604 3856
rect 287848 3816 287854 3828
rect 294598 3816 294604 3828
rect 294656 3816 294662 3868
rect 309042 3816 309048 3868
rect 309100 3856 309106 3868
rect 317322 3856 317328 3868
rect 309100 3828 317328 3856
rect 309100 3816 309106 3828
rect 317322 3816 317328 3828
rect 317380 3816 317386 3868
rect 330386 3816 330392 3868
rect 330444 3856 330450 3868
rect 341518 3856 341524 3868
rect 330444 3828 341524 3856
rect 330444 3816 330450 3828
rect 341518 3816 341524 3828
rect 341576 3816 341582 3868
rect 344554 3816 344560 3868
rect 344612 3856 344618 3868
rect 360838 3856 360844 3868
rect 344612 3828 360844 3856
rect 344612 3816 344618 3828
rect 360838 3816 360844 3828
rect 360896 3816 360902 3868
rect 365806 3816 365812 3868
rect 365864 3856 365870 3868
rect 400674 3856 400680 3868
rect 365864 3828 400680 3856
rect 365864 3816 365870 3828
rect 400674 3816 400680 3828
rect 400732 3816 400738 3868
rect 408402 3816 408408 3868
rect 408460 3856 408466 3868
rect 455414 3856 455420 3868
rect 408460 3828 455420 3856
rect 408460 3816 408466 3828
rect 455414 3816 455420 3828
rect 455472 3816 455478 3868
rect 495434 3816 495440 3868
rect 495492 3856 495498 3868
rect 564434 3856 564440 3868
rect 495492 3828 564440 3856
rect 495492 3816 495498 3828
rect 564434 3816 564440 3828
rect 564492 3816 564498 3868
rect 28902 3748 28908 3800
rect 28960 3788 28966 3800
rect 120074 3788 120080 3800
rect 28960 3760 120080 3788
rect 28960 3748 28966 3760
rect 120074 3748 120080 3760
rect 120132 3748 120138 3800
rect 142430 3748 142436 3800
rect 142488 3788 142494 3800
rect 305178 3788 305184 3800
rect 142488 3760 305184 3788
rect 142488 3748 142494 3760
rect 305178 3748 305184 3760
rect 305236 3748 305242 3800
rect 312630 3748 312636 3800
rect 312688 3788 312694 3800
rect 322198 3788 322204 3800
rect 312688 3760 322204 3788
rect 312688 3748 312694 3760
rect 322198 3748 322204 3760
rect 322256 3748 322262 3800
rect 323302 3748 323308 3800
rect 323360 3788 323366 3800
rect 335998 3788 336004 3800
rect 323360 3760 336004 3788
rect 323360 3748 323366 3760
rect 335998 3748 336004 3760
rect 336056 3748 336062 3800
rect 351638 3748 351644 3800
rect 351696 3788 351702 3800
rect 367830 3788 367836 3800
rect 351696 3760 367836 3788
rect 351696 3748 351702 3760
rect 367830 3748 367836 3760
rect 367888 3748 367894 3800
rect 369394 3748 369400 3800
rect 369452 3788 369458 3800
rect 403710 3788 403716 3800
rect 369452 3760 403716 3788
rect 369452 3748 369458 3760
rect 403710 3748 403716 3760
rect 403768 3748 403774 3800
rect 404814 3748 404820 3800
rect 404872 3788 404878 3800
rect 454218 3788 454224 3800
rect 404872 3760 454224 3788
rect 404872 3748 404878 3760
rect 454218 3748 454224 3760
rect 454276 3748 454282 3800
rect 496814 3748 496820 3800
rect 496872 3788 496878 3800
rect 568022 3788 568028 3800
rect 496872 3760 568028 3788
rect 496872 3748 496878 3760
rect 568022 3748 568028 3760
rect 568080 3748 568086 3800
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 118694 3720 118700 3732
rect 24268 3692 118700 3720
rect 24268 3680 24274 3692
rect 118694 3680 118700 3692
rect 118752 3680 118758 3732
rect 121086 3680 121092 3732
rect 121144 3720 121150 3732
rect 143626 3720 143632 3732
rect 121144 3692 143632 3720
rect 121144 3680 121150 3692
rect 143626 3680 143632 3692
rect 143684 3680 143690 3732
rect 145926 3680 145932 3732
rect 145984 3720 145990 3732
rect 356054 3720 356060 3732
rect 145984 3692 356060 3720
rect 145984 3680 145990 3692
rect 356054 3680 356060 3692
rect 356112 3680 356118 3732
rect 358722 3680 358728 3732
rect 358780 3720 358786 3732
rect 381538 3720 381544 3732
rect 358780 3692 381544 3720
rect 358780 3680 358786 3692
rect 381538 3680 381544 3692
rect 381596 3680 381602 3732
rect 387150 3680 387156 3732
rect 387208 3720 387214 3732
rect 448606 3720 448612 3732
rect 387208 3692 448612 3720
rect 387208 3680 387214 3692
rect 448606 3680 448612 3692
rect 448664 3680 448670 3732
rect 448698 3680 448704 3732
rect 448756 3720 448762 3732
rect 449802 3720 449808 3732
rect 448756 3692 449808 3720
rect 448756 3680 448762 3692
rect 449802 3680 449808 3692
rect 449860 3680 449866 3732
rect 496906 3680 496912 3732
rect 496964 3720 496970 3732
rect 571518 3720 571524 3732
rect 496964 3692 571524 3720
rect 496964 3680 496970 3692
rect 571518 3680 571524 3692
rect 571576 3680 571582 3732
rect 117590 3612 117596 3664
rect 117648 3652 117654 3664
rect 142154 3652 142160 3664
rect 117648 3624 142160 3652
rect 117648 3612 117654 3624
rect 142154 3612 142160 3624
rect 142212 3612 142218 3664
rect 147674 3652 147680 3664
rect 147646 3612 147680 3652
rect 147732 3612 147738 3664
rect 160186 3612 160192 3664
rect 160244 3652 160250 3664
rect 392118 3652 392124 3664
rect 160244 3624 392124 3652
rect 160244 3612 160250 3624
rect 392118 3612 392124 3624
rect 392176 3612 392182 3664
rect 401318 3612 401324 3664
rect 401376 3652 401382 3664
rect 454126 3652 454132 3664
rect 401376 3624 454132 3652
rect 401376 3612 401382 3624
rect 454126 3612 454132 3624
rect 454184 3612 454190 3664
rect 474918 3612 474924 3664
rect 474976 3652 474982 3664
rect 482830 3652 482836 3664
rect 474976 3624 482836 3652
rect 474976 3612 474982 3624
rect 482830 3612 482836 3624
rect 482888 3612 482894 3664
rect 498378 3612 498384 3664
rect 498436 3652 498442 3664
rect 575106 3652 575112 3664
rect 498436 3624 575112 3652
rect 498436 3612 498442 3624
rect 575106 3612 575112 3624
rect 575164 3612 575170 3664
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 147646 3584 147674 3612
rect 25372 3556 147674 3584
rect 25372 3544 25378 3556
rect 154206 3544 154212 3596
rect 154264 3584 154270 3596
rect 155218 3584 155224 3596
rect 154264 3556 155224 3584
rect 154264 3544 154270 3556
rect 155218 3544 155224 3556
rect 155276 3544 155282 3596
rect 156598 3544 156604 3596
rect 156656 3584 156662 3596
rect 390554 3584 390560 3596
rect 156656 3556 390560 3584
rect 156656 3544 156662 3556
rect 390554 3544 390560 3556
rect 390612 3544 390618 3596
rect 397730 3544 397736 3596
rect 397788 3584 397794 3596
rect 452654 3584 452660 3596
rect 397788 3556 452660 3584
rect 397788 3544 397794 3556
rect 452654 3544 452660 3556
rect 452712 3544 452718 3596
rect 464338 3544 464344 3596
rect 464396 3584 464402 3596
rect 474550 3584 474556 3596
rect 464396 3556 474556 3584
rect 464396 3544 464402 3556
rect 474550 3544 474556 3556
rect 474608 3544 474614 3596
rect 474826 3544 474832 3596
rect 474884 3584 474890 3596
rect 486418 3584 486424 3596
rect 474884 3556 486424 3584
rect 474884 3544 474890 3556
rect 486418 3544 486424 3556
rect 486476 3544 486482 3596
rect 499666 3544 499672 3596
rect 499724 3544 499730 3596
rect 502334 3544 502340 3596
rect 502392 3584 502398 3596
rect 582190 3584 582196 3596
rect 502392 3556 582196 3584
rect 502392 3544 502398 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 4798 3516 4804 3528
rect 1728 3488 4804 3516
rect 1728 3476 1734 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 20680 3488 147674 3516
rect 20680 3476 20686 3488
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 146386 3448 146392 3460
rect 15988 3420 146392 3448
rect 15988 3408 15994 3420
rect 146386 3408 146392 3420
rect 146444 3408 146450 3460
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 15838 3380 15844 3392
rect 11204 3352 15844 3380
rect 11204 3340 11210 3352
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 106918 3340 106924 3392
rect 106976 3380 106982 3392
rect 139394 3380 139400 3392
rect 106976 3352 139400 3380
rect 106976 3340 106982 3352
rect 139394 3340 139400 3352
rect 139452 3340 139458 3392
rect 147646 3380 147674 3488
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161290 3516 161296 3528
rect 160152 3488 161296 3516
rect 160152 3476 160158 3488
rect 161290 3476 161296 3488
rect 161348 3476 161354 3528
rect 161382 3476 161388 3528
rect 161440 3516 161446 3528
rect 389174 3516 389180 3528
rect 161440 3488 389180 3516
rect 161440 3476 161446 3488
rect 389174 3476 389180 3488
rect 389232 3476 389238 3528
rect 390646 3476 390652 3528
rect 390704 3516 390710 3528
rect 391842 3516 391848 3528
rect 390704 3488 391848 3516
rect 390704 3476 390710 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 398834 3476 398840 3528
rect 398892 3516 398898 3528
rect 400122 3516 400128 3528
rect 398892 3488 400128 3516
rect 398892 3476 398898 3488
rect 400122 3476 400128 3488
rect 400180 3476 400186 3528
rect 451366 3516 451372 3528
rect 400324 3488 451372 3516
rect 149514 3408 149520 3460
rect 149572 3448 149578 3460
rect 389266 3448 389272 3460
rect 149572 3420 389272 3448
rect 149572 3408 149578 3420
rect 389266 3408 389272 3420
rect 389324 3408 389330 3460
rect 390664 3420 393314 3448
rect 390664 3392 390692 3420
rect 147766 3380 147772 3392
rect 147646 3352 147772 3380
rect 147766 3340 147772 3352
rect 147824 3340 147830 3392
rect 153010 3340 153016 3392
rect 153068 3380 153074 3392
rect 161382 3380 161388 3392
rect 153068 3352 161388 3380
rect 153068 3340 153074 3352
rect 161382 3340 161388 3352
rect 161440 3340 161446 3392
rect 168374 3340 168380 3392
rect 168432 3380 168438 3392
rect 169570 3380 169576 3392
rect 168432 3352 169576 3380
rect 168432 3340 168438 3352
rect 169570 3340 169576 3352
rect 169628 3340 169634 3392
rect 201494 3340 201500 3392
rect 201552 3380 201558 3392
rect 202690 3380 202696 3392
rect 201552 3352 202696 3380
rect 201552 3340 201558 3352
rect 202690 3340 202696 3352
rect 202748 3340 202754 3392
rect 270034 3340 270040 3392
rect 270092 3380 270098 3392
rect 276658 3380 276664 3392
rect 270092 3352 276664 3380
rect 270092 3340 270098 3352
rect 276658 3340 276664 3352
rect 276716 3340 276722 3392
rect 299566 3340 299572 3392
rect 299624 3380 299630 3392
rect 300762 3380 300768 3392
rect 299624 3352 300768 3380
rect 299624 3340 299630 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 316126 3340 316132 3392
rect 316184 3380 316190 3392
rect 317322 3380 317328 3392
rect 316184 3352 317328 3380
rect 316184 3340 316190 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 390646 3340 390652 3392
rect 390704 3340 390710 3392
rect 110506 3272 110512 3324
rect 110564 3312 110570 3324
rect 140774 3312 140780 3324
rect 110564 3284 140780 3312
rect 110564 3272 110570 3284
rect 140774 3272 140780 3284
rect 140832 3272 140838 3324
rect 393286 3312 393314 3420
rect 394234 3340 394240 3392
rect 394292 3380 394298 3392
rect 400324 3380 400352 3488
rect 451366 3476 451372 3488
rect 451424 3476 451430 3528
rect 458082 3476 458088 3528
rect 458140 3516 458146 3528
rect 467926 3516 467932 3528
rect 458140 3488 467932 3516
rect 458140 3476 458146 3488
rect 467926 3476 467932 3488
rect 467984 3476 467990 3528
rect 476114 3476 476120 3528
rect 476172 3516 476178 3528
rect 489914 3516 489920 3528
rect 476172 3488 489920 3516
rect 476172 3476 476178 3488
rect 489914 3476 489920 3488
rect 489972 3476 489978 3528
rect 499684 3516 499712 3544
rect 578602 3516 578608 3528
rect 499684 3488 578608 3516
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 451274 3448 451280 3460
rect 394292 3352 400352 3380
rect 402946 3420 451280 3448
rect 394292 3340 394298 3352
rect 402946 3312 402974 3420
rect 451274 3408 451280 3420
rect 451332 3408 451338 3460
rect 461670 3408 461676 3460
rect 461728 3448 461734 3460
rect 478138 3448 478144 3460
rect 461728 3420 478144 3448
rect 461728 3408 461734 3420
rect 478138 3408 478144 3420
rect 478196 3408 478202 3460
rect 500954 3408 500960 3460
rect 501012 3448 501018 3460
rect 580994 3448 581000 3460
rect 501012 3420 581000 3448
rect 501012 3408 501018 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 426158 3340 426164 3392
rect 426216 3380 426222 3392
rect 459554 3380 459560 3392
rect 426216 3352 459560 3380
rect 426216 3340 426222 3352
rect 459554 3340 459560 3352
rect 459612 3340 459618 3392
rect 491386 3340 491392 3392
rect 491444 3380 491450 3392
rect 546678 3380 546684 3392
rect 491444 3352 546684 3380
rect 491444 3340 491450 3352
rect 546678 3340 546684 3352
rect 546736 3340 546742 3392
rect 393286 3284 402974 3312
rect 433242 3272 433248 3324
rect 433300 3312 433306 3324
rect 462498 3312 462504 3324
rect 433300 3284 462504 3312
rect 433300 3272 433306 3284
rect 462498 3272 462504 3284
rect 462556 3272 462562 3324
rect 490006 3272 490012 3324
rect 490064 3312 490070 3324
rect 543182 3312 543188 3324
rect 490064 3284 543188 3312
rect 490064 3272 490070 3284
rect 543182 3272 543188 3284
rect 543240 3272 543246 3324
rect 13538 3204 13544 3256
rect 13596 3244 13602 3256
rect 14458 3244 14464 3256
rect 13596 3216 14464 3244
rect 13596 3204 13602 3216
rect 14458 3204 14464 3216
rect 14516 3204 14522 3256
rect 114002 3204 114008 3256
rect 114060 3244 114066 3256
rect 142246 3244 142252 3256
rect 114060 3216 142252 3244
rect 114060 3204 114066 3216
rect 142246 3204 142252 3216
rect 142304 3204 142310 3256
rect 440326 3204 440332 3256
rect 440384 3244 440390 3256
rect 441522 3244 441528 3256
rect 440384 3216 441528 3244
rect 440384 3204 440390 3216
rect 441522 3204 441528 3216
rect 441580 3204 441586 3256
rect 443822 3204 443828 3256
rect 443880 3244 443886 3256
rect 465074 3244 465080 3256
rect 443880 3216 465080 3244
rect 443880 3204 443886 3216
rect 465074 3204 465080 3216
rect 465132 3204 465138 3256
rect 488534 3204 488540 3256
rect 488592 3244 488598 3256
rect 539594 3244 539600 3256
rect 488592 3216 539600 3244
rect 488592 3204 488598 3216
rect 539594 3204 539600 3216
rect 539652 3204 539658 3256
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 117498 3176 117504 3188
rect 19484 3148 117504 3176
rect 19484 3136 19490 3148
rect 117498 3136 117504 3148
rect 117556 3136 117562 3188
rect 280706 3136 280712 3188
rect 280764 3176 280770 3188
rect 284938 3176 284944 3188
rect 280764 3148 284944 3176
rect 280764 3136 280770 3148
rect 284938 3136 284944 3148
rect 284996 3136 285002 3188
rect 531314 3136 531320 3188
rect 531372 3176 531378 3188
rect 532142 3176 532148 3188
rect 531372 3148 532148 3176
rect 531372 3136 531378 3148
rect 532142 3136 532148 3148
rect 532200 3136 532206 3188
rect 316034 3068 316040 3120
rect 316092 3108 316098 3120
rect 318518 3108 318524 3120
rect 316092 3080 318524 3108
rect 316092 3068 316098 3080
rect 318518 3068 318524 3080
rect 318576 3068 318582 3120
rect 316218 3000 316224 3052
rect 316276 3040 316282 3052
rect 324958 3040 324964 3052
rect 316276 3012 324964 3040
rect 316276 3000 316282 3012
rect 324958 3000 324964 3012
rect 325016 3000 325022 3052
rect 473354 3000 473360 3052
rect 473412 3040 473418 3052
rect 479334 3040 479340 3052
rect 473412 3012 479340 3040
rect 473412 3000 473418 3012
rect 479334 3000 479340 3012
rect 479392 3000 479398 3052
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 11698 2972 11704 2984
rect 10008 2944 11704 2972
rect 10008 2932 10014 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 298462 2864 298468 2916
rect 298520 2904 298526 2916
rect 304258 2904 304264 2916
rect 298520 2876 304264 2904
rect 298520 2864 298526 2876
rect 304258 2864 304264 2876
rect 304316 2864 304322 2916
rect 199102 2320 199108 2372
rect 199160 2360 199166 2372
rect 401594 2360 401600 2372
rect 199160 2332 401600 2360
rect 199160 2320 199166 2332
rect 401594 2320 401600 2332
rect 401652 2320 401658 2372
rect 192018 2252 192024 2304
rect 192076 2292 192082 2304
rect 400398 2292 400404 2304
rect 192076 2264 400404 2292
rect 192076 2252 192082 2264
rect 400398 2252 400404 2264
rect 400456 2252 400462 2304
rect 181438 2184 181444 2236
rect 181496 2224 181502 2236
rect 396718 2224 396724 2236
rect 181496 2196 396724 2224
rect 181496 2184 181502 2196
rect 396718 2184 396724 2196
rect 396776 2184 396782 2236
rect 167178 2116 167184 2168
rect 167236 2156 167242 2168
rect 393314 2156 393320 2168
rect 167236 2128 393320 2156
rect 167236 2116 167242 2128
rect 393314 2116 393320 2128
rect 393372 2116 393378 2168
rect 237374 2048 237380 2100
rect 237432 2088 237438 2100
rect 466270 2088 466276 2100
rect 237432 2060 466276 2088
rect 237432 2048 237438 2060
rect 466270 2048 466276 2060
rect 466328 2048 466334 2100
<< via1 >>
rect 56600 29860 56652 29912
rect 57643 29860 57695 29912
rect 62120 29860 62172 29912
rect 63100 29860 63152 29912
rect 71872 29792 71924 29844
rect 73079 29792 73131 29844
rect 77300 29792 77352 29844
rect 78553 29792 78605 29844
rect 80060 29792 80112 29844
rect 81290 29792 81342 29844
rect 82820 29792 82872 29844
rect 83993 29792 84045 29844
rect 85672 29792 85724 29844
rect 86730 29792 86782 29844
rect 88432 29792 88484 29844
rect 89450 29792 89502 29844
rect 111892 29792 111944 29844
rect 113097 29792 113149 29844
rect 128360 29792 128412 29844
rect 129485 29792 129537 29844
rect 133880 29792 133932 29844
rect 134942 29792 134994 29844
rect 136640 29792 136692 29844
rect 137679 29792 137731 29844
rect 139400 29792 139452 29844
rect 140399 29792 140451 29844
rect 189080 29792 189132 29844
rect 190413 29792 190465 29844
rect 197452 29792 197504 29844
rect 198573 29792 198625 29844
rect 200120 29792 200172 29844
rect 201310 29792 201362 29844
rect 205640 29792 205692 29844
rect 206750 29792 206802 29844
rect 211160 29792 211212 29844
rect 212241 29792 212293 29844
rect 231860 29792 231912 29844
rect 233134 29792 233186 29844
rect 237380 29792 237432 29844
rect 238608 29792 238660 29844
rect 240140 29792 240192 29844
rect 241362 29792 241414 29844
rect 242900 29792 242952 29844
rect 244048 29792 244100 29844
rect 259460 29792 259512 29844
rect 260436 29792 260488 29844
rect 274640 29792 274692 29844
rect 275889 29792 275941 29844
rect 277492 29792 277544 29844
rect 278609 29792 278661 29844
rect 285680 29792 285732 29844
rect 286837 29792 286889 29844
rect 291200 29792 291252 29844
rect 292260 29792 292312 29844
rect 311900 29792 311952 29844
rect 313153 29792 313205 29844
rect 314752 29792 314804 29844
rect 315890 29792 315942 29844
rect 317420 29792 317472 29844
rect 318627 29792 318679 29844
rect 346400 29792 346452 29844
rect 347731 29792 347783 29844
rect 352012 29792 352064 29844
rect 353188 29792 353240 29844
rect 357440 29792 357492 29844
rect 358645 29792 358697 29844
rect 362960 29792 363012 29844
rect 364102 29792 364154 29844
rect 374000 29792 374052 29844
rect 375016 29792 375068 29844
rect 389180 29792 389232 29844
rect 390469 29792 390521 29844
rect 405740 29792 405792 29844
rect 406857 29792 406909 29844
rect 426532 29792 426584 29844
rect 427750 29792 427802 29844
rect 431960 29792 432012 29844
rect 433173 29792 433225 29844
rect 434812 29792 434864 29844
rect 435927 29792 435979 29844
rect 448520 29792 448572 29844
rect 449578 29792 449630 29844
rect 474832 29792 474884 29844
rect 475979 29792 476031 29844
rect 488540 29792 488592 29844
rect 489613 29792 489665 29844
rect 491300 29792 491352 29844
rect 492316 29792 492368 29844
rect 494060 29792 494112 29844
rect 495053 29792 495105 29844
rect 201500 28500 201552 28552
rect 403164 28500 403216 28552
rect 194600 28432 194652 28484
rect 401416 28432 401468 28484
rect 185032 28364 185084 28416
rect 398656 28364 398708 28416
rect 176660 28296 176712 28348
rect 396816 28296 396868 28348
rect 162860 28228 162912 28280
rect 393228 28228 393280 28280
rect 64880 28092 64932 28144
rect 65800 28092 65852 28144
rect 67640 28092 67692 28144
rect 68560 28092 68612 28144
rect 102140 28092 102192 28144
rect 103060 28092 103112 28144
rect 104900 28092 104952 28144
rect 105820 28092 105872 28144
rect 110420 28092 110472 28144
rect 111248 28092 111300 28144
rect 114652 28092 114704 28144
rect 115848 28092 115900 28144
rect 142160 28092 142212 28144
rect 143080 28092 143132 28144
rect 147680 28092 147732 28144
rect 148508 28092 148560 28144
rect 151912 28092 151964 28144
rect 153108 28092 153160 28144
rect 182180 28092 182232 28144
rect 183100 28092 183152 28144
rect 222200 28092 222252 28144
rect 223120 28092 223172 28144
rect 269212 28092 269264 28144
rect 270408 28092 270460 28144
rect 302240 28092 302292 28144
rect 303160 28092 303212 28144
rect 309232 28092 309284 28144
rect 310428 28092 310480 28144
rect 339500 28092 339552 28144
rect 340420 28092 340472 28144
rect 429292 28092 429344 28144
rect 430488 28092 430540 28144
rect 456800 28092 456852 28144
rect 457720 28092 457772 28144
rect 459560 28092 459612 28144
rect 460480 28092 460532 28144
rect 69020 27548 69072 27600
rect 72148 27548 72200 27600
rect 90364 27548 90416 27600
rect 92204 27548 92256 27600
rect 106924 27548 106976 27600
rect 107660 27548 107712 27600
rect 108948 27548 109000 27600
rect 109500 27548 109552 27600
rect 114008 27548 114060 27600
rect 115940 27548 115992 27600
rect 117228 27548 117280 27600
rect 117688 27548 117740 27600
rect 126244 27548 126296 27600
rect 127624 27548 127676 27600
rect 155224 27548 155276 27600
rect 158536 27548 158588 27600
rect 163136 27548 163188 27600
rect 170404 27548 170456 27600
rect 171324 27548 171376 27600
rect 173164 27548 173216 27600
rect 185860 27548 185912 27600
rect 186964 27548 187016 27600
rect 204076 27548 204128 27600
rect 205548 27548 205600 27600
rect 243176 27548 243228 27600
rect 244924 27548 244976 27600
rect 254032 27548 254084 27600
rect 256608 27548 256660 27600
rect 264980 27548 265032 27600
rect 267648 27548 267700 27600
rect 282184 27548 282236 27600
rect 283196 27548 283248 27600
rect 300124 27548 300176 27600
rect 301320 27548 301372 27600
rect 313924 27548 313976 27600
rect 314936 27548 314988 27600
rect 325884 27548 325936 27600
rect 327724 27548 327776 27600
rect 355968 27548 356020 27600
rect 356704 27548 356756 27600
rect 396724 27548 396776 27600
rect 397736 27548 397788 27600
rect 407764 27548 407816 27600
rect 408684 27548 408736 27600
rect 416688 27548 416740 27600
rect 421288 27548 421340 27600
rect 425704 27548 425756 27600
rect 428648 27548 428700 27600
rect 465264 27548 465316 27600
rect 470508 27548 470560 27600
rect 473268 27548 473320 27600
rect 474740 27548 474792 27600
rect 481364 27548 481416 27600
rect 485044 27548 485096 27600
rect 109040 27480 109092 27532
rect 112168 27480 112220 27532
rect 225880 27480 225932 27532
rect 249064 27480 249116 27532
rect 298744 27480 298796 27532
rect 300400 27480 300452 27532
rect 361396 27480 361448 27532
rect 376116 27480 376168 27532
rect 461032 27480 461084 27532
rect 469588 27480 469640 27532
rect 214932 27412 214984 27464
rect 273904 27412 273956 27464
rect 368664 27412 368716 27464
rect 414664 27412 414716 27464
rect 207664 27344 207716 27396
rect 291844 27344 291896 27396
rect 336832 27344 336884 27396
rect 353392 27344 353444 27396
rect 362316 27344 362368 27396
rect 410524 27344 410576 27396
rect 413284 27344 413336 27396
rect 426808 27344 426860 27396
rect 203156 27276 203208 27328
rect 296076 27276 296128 27328
rect 348608 27276 348660 27328
rect 364984 27276 365036 27328
rect 367744 27276 367796 27328
rect 419540 27276 419592 27328
rect 454040 27276 454092 27328
rect 467748 27276 467800 27328
rect 95148 27208 95200 27260
rect 95792 27208 95844 27260
rect 219532 27208 219584 27260
rect 339132 27208 339184 27260
rect 341340 27208 341392 27260
rect 360476 27208 360528 27260
rect 380440 27208 380492 27260
rect 453304 27208 453356 27260
rect 130384 27140 130436 27192
rect 131304 27140 131356 27192
rect 196808 27140 196860 27192
rect 242164 27140 242216 27192
rect 261392 27140 261444 27192
rect 407856 27140 407908 27192
rect 410432 27140 410484 27192
rect 415952 27140 416004 27192
rect 418804 27140 418856 27192
rect 440424 27140 440476 27192
rect 449900 27140 449952 27192
rect 466828 27140 466880 27192
rect 184940 27072 184992 27124
rect 246304 27072 246356 27124
rect 249524 27072 249576 27124
rect 396816 27072 396868 27124
rect 403624 27072 403676 27124
rect 437756 27072 437808 27124
rect 447232 27072 447284 27124
rect 466000 27072 466052 27124
rect 480444 27072 480496 27124
rect 503720 27072 503772 27124
rect 143540 27004 143592 27056
rect 155868 27004 155920 27056
rect 166816 27004 166868 27056
rect 184204 27004 184256 27056
rect 189448 27004 189500 27056
rect 199384 27004 199436 27056
rect 240416 27004 240468 27056
rect 418896 27004 418948 27056
rect 421564 27004 421616 27056
rect 425888 27004 425940 27056
rect 440240 27004 440292 27056
rect 464160 27004 464212 27056
rect 485964 27004 486016 27056
rect 512644 27004 512696 27056
rect 15844 26936 15896 26988
rect 145840 26936 145892 26988
rect 146300 26936 146352 26988
rect 156788 26936 156840 26988
rect 172244 26936 172296 26988
rect 191104 26936 191156 26988
rect 191932 26936 191984 26988
rect 193128 26936 193180 26988
rect 242256 26936 242308 26988
rect 424324 26936 424376 26988
rect 424416 26936 424468 26988
rect 434996 26936 435048 26988
rect 436100 26936 436152 26988
rect 463240 26936 463292 26988
rect 482284 26936 482336 26988
rect 510620 26936 510672 26988
rect 10324 26868 10376 26920
rect 149520 26868 149572 26920
rect 150440 26868 150492 26920
rect 157708 26868 157760 26920
rect 161296 26868 161348 26920
rect 164240 26868 164292 26920
rect 167644 26868 167696 26920
rect 175924 26868 175976 26920
rect 176752 26868 176804 26920
rect 224224 26868 224276 26920
rect 230388 26868 230440 26920
rect 428464 26868 428516 26920
rect 429384 26868 429436 26920
rect 461400 26868 461452 26920
rect 477776 26868 477828 26920
rect 492680 26868 492732 26920
rect 500500 26868 500552 26920
rect 569224 26868 569276 26920
rect 271972 26800 272024 26852
rect 273168 26800 273220 26852
rect 157524 26664 157576 26716
rect 159456 26664 159508 26716
rect 77668 26324 77720 26376
rect 79324 26324 79376 26376
rect 93124 26324 93176 26376
rect 94044 26324 94096 26376
rect 54484 26256 54536 26308
rect 55864 26256 55916 26308
rect 74080 26256 74132 26308
rect 75920 26256 75972 26308
rect 295984 26256 296036 26308
rect 296812 26324 296864 26376
rect 379612 26324 379664 26376
rect 381544 26324 381596 26376
rect 421012 26256 421064 26308
rect 424048 26256 424100 26308
rect 467840 26256 467892 26308
rect 471336 26256 471388 26308
rect 478696 26256 478748 26308
rect 482284 26256 482336 26308
rect 382280 26188 382332 26240
rect 383200 26188 383252 26240
rect 386420 26188 386472 26240
rect 387708 26188 387760 26240
rect 353392 26120 353444 26172
rect 396080 26120 396132 26172
rect 70400 26052 70452 26104
rect 71228 26052 71280 26104
rect 74632 26052 74684 26104
rect 75828 26052 75880 26104
rect 376024 26052 376076 26104
rect 441620 26052 441672 26104
rect 200212 25984 200264 26036
rect 316132 25984 316184 26036
rect 343640 25984 343692 26036
rect 423680 25984 423732 26036
rect 197360 25916 197412 25968
rect 285772 25916 285824 25968
rect 312544 25916 312596 25968
rect 429200 25916 429252 25968
rect 208492 25848 208544 25900
rect 351920 25848 351972 25900
rect 356060 25848 356112 25900
rect 464344 25848 464396 25900
rect 216772 25780 216824 25832
rect 383660 25780 383712 25832
rect 231952 25712 232004 25764
rect 440332 25712 440384 25764
rect 84200 25644 84252 25696
rect 118792 25644 118844 25696
rect 247040 25644 247092 25696
rect 501052 25644 501104 25696
rect 4804 25576 4856 25628
rect 55312 25576 55364 25628
rect 88340 25576 88392 25628
rect 135260 25576 135312 25628
rect 259552 25576 259604 25628
rect 547880 25576 547932 25628
rect 27620 25508 27672 25560
rect 91008 25508 91060 25560
rect 183560 25508 183612 25560
rect 252560 25508 252612 25560
rect 266360 25508 266412 25560
rect 575480 25508 575532 25560
rect 345112 24692 345164 24744
rect 432144 24692 432196 24744
rect 189080 24624 189132 24676
rect 277400 24624 277452 24676
rect 339132 24624 339184 24676
rect 390652 24624 390704 24676
rect 198740 24556 198792 24608
rect 313280 24556 313332 24608
rect 330484 24556 330536 24608
rect 431960 24556 432012 24608
rect 276664 24488 276716 24540
rect 419632 24488 419684 24540
rect 205732 24420 205784 24472
rect 338120 24420 338172 24472
rect 367100 24420 367152 24472
rect 516140 24420 516192 24472
rect 213920 24352 213972 24404
rect 369860 24352 369912 24404
rect 385684 24352 385736 24404
rect 447140 24352 447192 24404
rect 224960 24284 225012 24336
rect 412640 24284 412692 24336
rect 46940 24216 46992 24268
rect 66260 24216 66312 24268
rect 69112 24216 69164 24268
rect 102232 24216 102284 24268
rect 236000 24216 236052 24268
rect 458272 24216 458324 24268
rect 44180 24148 44232 24200
rect 95148 24148 95200 24200
rect 99380 24148 99432 24200
rect 138020 24148 138072 24200
rect 248420 24148 248472 24200
rect 505100 24148 505152 24200
rect 13820 24080 13872 24132
rect 117228 24080 117280 24132
rect 176752 24080 176804 24132
rect 227720 24080 227772 24132
rect 259460 24080 259512 24132
rect 550640 24080 550692 24132
rect 336740 23332 336792 23384
rect 398840 23332 398892 23384
rect 197544 23264 197596 23316
rect 306472 23264 306524 23316
rect 341524 23264 341576 23316
rect 434812 23264 434864 23316
rect 205640 23196 205692 23248
rect 340880 23196 340932 23248
rect 354680 23196 354732 23248
rect 466460 23196 466512 23248
rect 147864 23128 147916 23180
rect 271972 23128 272024 23180
rect 273260 23128 273312 23180
rect 416688 23128 416740 23180
rect 215300 23060 215352 23112
rect 376760 23060 376812 23112
rect 129832 22992 129884 23044
rect 267832 22992 267884 23044
rect 371332 22992 371384 23044
rect 534080 22992 534132 23044
rect 51080 22924 51132 22976
rect 67732 22924 67784 22976
rect 227904 22924 227956 22976
rect 426440 22924 426492 22976
rect 87052 22856 87104 22908
rect 106280 22856 106332 22908
rect 245752 22856 245804 22908
rect 498292 22856 498344 22908
rect 67732 22788 67784 22840
rect 129740 22788 129792 22840
rect 253940 22788 253992 22840
rect 529940 22788 529992 22840
rect 22100 22720 22152 22772
rect 89720 22720 89772 22772
rect 173992 22720 174044 22772
rect 218060 22720 218112 22772
rect 264980 22720 265032 22772
rect 572720 22720 572772 22772
rect 193312 21972 193364 22024
rect 284300 21972 284352 22024
rect 367836 21972 367888 22024
rect 440424 21972 440476 22024
rect 197452 21904 197504 21956
rect 309324 21904 309376 21956
rect 342352 21904 342404 21956
rect 420920 21904 420972 21956
rect 143724 21836 143776 21888
rect 271880 21836 271932 21888
rect 322204 21836 322256 21888
rect 430580 21836 430632 21888
rect 251180 21768 251232 21820
rect 410432 21768 410484 21820
rect 216680 21700 216732 21752
rect 380992 21700 381044 21752
rect 208400 21632 208452 21684
rect 349160 21632 349212 21684
rect 372620 21632 372672 21684
rect 538220 21632 538272 21684
rect 229100 21564 229152 21616
rect 430580 21564 430632 21616
rect 80152 21496 80204 21548
rect 104992 21496 105044 21548
rect 244280 21496 244332 21548
rect 490012 21496 490064 21548
rect 16580 21428 16632 21480
rect 59268 21428 59320 21480
rect 74724 21428 74776 21480
rect 131212 21428 131264 21480
rect 252652 21428 252704 21480
rect 523040 21428 523092 21480
rect 34520 21360 34572 21412
rect 92480 21360 92532 21412
rect 173900 21360 173952 21412
rect 213920 21360 213972 21412
rect 263600 21360 263652 21412
rect 564532 21360 564584 21412
rect 360476 20544 360528 20596
rect 414204 20544 414256 20596
rect 325700 20476 325752 20528
rect 424416 20476 424468 20528
rect 205548 20408 205600 20460
rect 331404 20408 331456 20460
rect 346492 20408 346544 20460
rect 434720 20408 434772 20460
rect 136824 20340 136876 20392
rect 269212 20340 269264 20392
rect 284300 20340 284352 20392
rect 421012 20340 421064 20392
rect 211160 20272 211212 20324
rect 363144 20272 363196 20324
rect 219440 20204 219492 20256
rect 394884 20204 394936 20256
rect 20720 20136 20772 20188
rect 59452 20136 59504 20188
rect 234712 20136 234764 20188
rect 455512 20136 455564 20188
rect 98092 20068 98144 20120
rect 108948 20068 109000 20120
rect 245660 20068 245712 20120
rect 494244 20068 494296 20120
rect 59360 20000 59412 20052
rect 99288 20000 99340 20052
rect 172520 20000 172572 20052
rect 209872 20000 209924 20052
rect 256608 20000 256660 20052
rect 525800 20000 525852 20052
rect 52460 19932 52512 19984
rect 125692 19932 125744 19984
rect 186320 19932 186372 19984
rect 263600 19932 263652 19984
rect 267648 19932 267700 19984
rect 568580 19932 568632 19984
rect 342260 19184 342312 19236
rect 416964 19184 417016 19236
rect 364984 19116 365036 19168
rect 441620 19116 441672 19168
rect 140872 19048 140924 19100
rect 270500 19048 270552 19100
rect 304264 19048 304316 19100
rect 426532 19048 426584 19100
rect 204260 18980 204312 19032
rect 334164 18980 334216 19032
rect 353944 18980 353996 19032
rect 437572 18980 437624 19032
rect 212540 18912 212592 18964
rect 365904 18912 365956 18964
rect 29000 18844 29052 18896
rect 62212 18844 62264 18896
rect 220820 18844 220872 18896
rect 398932 18844 398984 18896
rect 237472 18776 237524 18828
rect 462412 18776 462464 18828
rect 62212 18708 62264 18760
rect 99472 18708 99524 18760
rect 242900 18708 242952 18760
rect 487160 18708 487212 18760
rect 487252 18708 487304 18760
rect 531320 18708 531372 18760
rect 92480 18640 92532 18692
rect 136732 18640 136784 18692
rect 169760 18640 169812 18692
rect 200212 18640 200264 18692
rect 251364 18640 251416 18692
rect 518900 18640 518952 18692
rect 49700 18572 49752 18624
rect 125600 18572 125652 18624
rect 186964 18572 187016 18624
rect 259460 18572 259512 18624
rect 262312 18572 262364 18624
rect 561680 18572 561732 18624
rect 211160 17756 211212 17808
rect 288532 17756 288584 17808
rect 345020 17756 345072 17808
rect 427820 17756 427872 17808
rect 201592 17688 201644 17740
rect 324412 17688 324464 17740
rect 324964 17688 325016 17740
rect 432052 17688 432104 17740
rect 211252 17620 211304 17672
rect 358912 17620 358964 17672
rect 374092 17620 374144 17672
rect 540980 17620 541032 17672
rect 218152 17552 218204 17604
rect 387892 17552 387944 17604
rect 226432 17484 226484 17536
rect 408592 17484 408644 17536
rect 233240 17416 233292 17468
rect 448796 17416 448848 17468
rect 73160 17348 73212 17400
rect 102140 17348 102192 17400
rect 244924 17348 244976 17400
rect 483204 17348 483256 17400
rect 35900 17280 35952 17332
rect 63500 17280 63552 17332
rect 81532 17280 81584 17332
rect 133972 17280 134024 17332
rect 168472 17280 168524 17332
rect 195980 17280 196032 17332
rect 251272 17280 251324 17332
rect 514760 17280 514812 17332
rect 41420 17212 41472 17264
rect 93952 17212 94004 17264
rect 180800 17212 180852 17264
rect 242900 17212 242952 17264
rect 262220 17212 262272 17264
rect 557540 17212 557592 17264
rect 411904 16532 411956 16584
rect 448612 16532 448664 16584
rect 208584 16464 208636 16516
rect 288440 16464 288492 16516
rect 342904 16464 342956 16516
rect 436192 16464 436244 16516
rect 183744 16396 183796 16448
rect 281540 16396 281592 16448
rect 357532 16396 357584 16448
rect 461676 16396 461728 16448
rect 259552 16328 259604 16380
rect 416872 16328 416924 16380
rect 255872 16260 255924 16312
rect 416780 16260 416832 16312
rect 248420 16192 248472 16244
rect 414112 16192 414164 16244
rect 245200 16124 245252 16176
rect 414020 16124 414072 16176
rect 126980 16056 127032 16108
rect 267740 16056 267792 16108
rect 374000 16056 374052 16108
rect 545488 16056 545540 16108
rect 241704 15988 241756 16040
rect 412732 15988 412784 16040
rect 40224 15920 40276 15972
rect 64972 15920 65024 15972
rect 66720 15920 66772 15972
rect 100760 15920 100812 15972
rect 102232 15920 102284 15972
rect 110512 15920 110564 15972
rect 132960 15920 133012 15972
rect 151912 15920 151964 15972
rect 168380 15920 168432 15972
rect 193404 15920 193456 15972
rect 237656 15920 237708 15972
rect 411352 15920 411404 15972
rect 418896 15920 418948 15972
rect 473452 15920 473504 15972
rect 488632 15920 488684 15972
rect 536104 15920 536156 15972
rect 11704 15852 11756 15904
rect 116032 15852 116084 15904
rect 138848 15852 138900 15904
rect 386512 15852 386564 15904
rect 414664 15852 414716 15904
rect 520280 15852 520332 15904
rect 378784 15104 378836 15156
rect 443092 15104 443144 15156
rect 336004 15036 336056 15088
rect 433340 15036 433392 15088
rect 294604 14968 294656 15020
rect 425152 14968 425204 15020
rect 231032 14900 231084 14952
rect 409880 14900 409932 14952
rect 381544 14832 381596 14884
rect 563060 14832 563112 14884
rect 219992 14764 220044 14816
rect 407120 14764 407172 14816
rect 216864 14696 216916 14748
rect 405740 14696 405792 14748
rect 213368 14628 213420 14680
rect 405832 14628 405884 14680
rect 82912 14560 82964 14612
rect 111616 14560 111668 14612
rect 209964 14560 210016 14612
rect 404360 14560 404412 14612
rect 405004 14560 405056 14612
rect 445852 14560 445904 14612
rect 60832 14492 60884 14544
rect 128452 14492 128504 14544
rect 206192 14492 206244 14544
rect 403072 14492 403124 14544
rect 410524 14492 410576 14544
rect 495532 14492 495584 14544
rect 14464 14424 14516 14476
rect 88524 14424 88576 14476
rect 135260 14424 135312 14476
rect 385132 14424 385184 14476
rect 407856 14424 407908 14476
rect 554780 14424 554832 14476
rect 268384 13676 268436 13728
rect 303620 13676 303672 13728
rect 346400 13676 346452 13728
rect 439136 13676 439188 13728
rect 273904 13608 273956 13660
rect 374092 13608 374144 13660
rect 158904 13540 158956 13592
rect 274640 13540 274692 13592
rect 376116 13540 376168 13592
rect 492312 13540 492364 13592
rect 154672 13472 154724 13524
rect 274732 13472 274784 13524
rect 284944 13472 284996 13524
rect 422392 13472 422444 13524
rect 152004 13404 152056 13456
rect 273352 13404 273404 13456
rect 369952 13404 370004 13456
rect 527824 13404 527876 13456
rect 249064 13336 249116 13388
rect 415400 13336 415452 13388
rect 234620 13268 234672 13320
rect 451648 13268 451700 13320
rect 80244 13200 80296 13252
rect 100760 13200 100812 13252
rect 173900 13200 173952 13252
rect 394792 13200 394844 13252
rect 64328 13132 64380 13184
rect 128360 13132 128412 13184
rect 170312 13132 170364 13184
rect 394700 13132 394752 13184
rect 485780 13132 485832 13184
rect 528560 13132 528612 13184
rect 17960 13064 18012 13116
rect 88432 13064 88484 13116
rect 128176 13064 128228 13116
rect 383752 13064 383804 13116
rect 396816 13064 396868 13116
rect 508872 13064 508924 13116
rect 360844 12996 360896 13048
rect 438860 12996 438912 13048
rect 105728 12452 105780 12504
rect 110420 12452 110472 12504
rect 327724 12384 327776 12436
rect 353576 12384 353628 12436
rect 261760 12316 261812 12368
rect 302332 12316 302384 12368
rect 325792 12316 325844 12368
rect 357532 12316 357584 12368
rect 247592 12248 247644 12300
rect 298100 12248 298152 12300
rect 349252 12248 349304 12300
rect 445852 12248 445904 12300
rect 236552 12180 236604 12232
rect 295340 12180 295392 12232
rect 349344 12180 349396 12232
rect 448704 12180 448756 12232
rect 233424 12112 233476 12164
rect 294052 12112 294104 12164
rect 350540 12112 350592 12164
rect 453304 12112 453356 12164
rect 226524 12044 226576 12096
rect 292580 12044 292632 12096
rect 299572 12044 299624 12096
rect 311992 12044 312044 12096
rect 352104 12044 352156 12096
rect 457076 12044 457128 12096
rect 222752 11976 222804 12028
rect 291200 11976 291252 12028
rect 296076 11976 296128 12028
rect 328000 11976 328052 12028
rect 352012 11976 352064 12028
rect 459928 11976 459980 12028
rect 77300 11908 77352 11960
rect 93952 11908 94004 11960
rect 219256 11908 219308 11960
rect 291292 11908 291344 11960
rect 291844 11908 291896 11960
rect 345296 11908 345348 11960
rect 353300 11908 353352 11960
rect 463976 11908 464028 11960
rect 84200 11840 84252 11892
rect 104900 11840 104952 11892
rect 215300 11840 215352 11892
rect 289820 11840 289872 11892
rect 294512 11840 294564 11892
rect 413284 11840 413336 11892
rect 485044 11840 485096 11892
rect 507216 11840 507268 11892
rect 44272 11772 44324 11824
rect 64880 11772 64932 11824
rect 85764 11772 85816 11824
rect 133880 11772 133932 11824
rect 133972 11772 134024 11824
rect 269120 11772 269172 11824
rect 273904 11772 273956 11824
rect 418160 11772 418212 11824
rect 484400 11772 484452 11824
rect 521660 11772 521712 11824
rect 30840 11704 30892 11756
rect 90364 11704 90416 11756
rect 188528 11704 188580 11756
rect 399024 11704 399076 11756
rect 453396 11704 453448 11756
rect 566832 11704 566884 11756
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 264980 10956 265032 11008
rect 302240 10956 302292 11008
rect 311440 10956 311492 11008
rect 313924 10956 313976 11008
rect 334072 10956 334124 11008
rect 389456 10956 389508 11008
rect 251272 10888 251324 10940
rect 299664 10888 299716 10940
rect 335360 10888 335412 10940
rect 392032 10888 392084 10940
rect 229376 10820 229428 10872
rect 293960 10820 294012 10872
rect 381544 10820 381596 10872
rect 443000 10820 443052 10872
rect 180248 10752 180300 10804
rect 280252 10752 280304 10804
rect 338212 10752 338264 10804
rect 403532 10752 403584 10804
rect 403716 10752 403768 10804
rect 445760 10752 445812 10804
rect 172704 10684 172756 10736
rect 278780 10684 278832 10736
rect 339592 10684 339644 10736
rect 407212 10684 407264 10736
rect 168380 10616 168432 10668
rect 277492 10616 277544 10668
rect 339500 10616 339552 10668
rect 410800 10616 410852 10668
rect 166080 10548 166132 10600
rect 277584 10548 277636 10600
rect 301504 10548 301556 10600
rect 425704 10548 425756 10600
rect 269764 10480 269816 10532
rect 411260 10480 411312 10532
rect 77392 10412 77444 10464
rect 103520 10412 103572 10464
rect 162032 10412 162084 10464
rect 276020 10412 276072 10464
rect 283104 10412 283156 10464
rect 306564 10412 306616 10464
rect 371240 10412 371292 10464
rect 531412 10412 531464 10464
rect 33600 10344 33652 10396
rect 62120 10344 62172 10396
rect 78680 10344 78732 10396
rect 97448 10344 97500 10396
rect 103336 10344 103388 10396
rect 139492 10344 139544 10396
rect 238760 10344 238812 10396
rect 469864 10344 469916 10396
rect 478880 10344 478932 10396
rect 499580 10344 499632 10396
rect 56784 10276 56836 10328
rect 126244 10276 126296 10328
rect 240140 10276 240192 10328
rect 476488 10276 476540 10328
rect 483112 10276 483164 10328
rect 517888 10276 517940 10328
rect 400680 9528 400732 9580
rect 444380 9528 444432 9580
rect 254676 9460 254728 9512
rect 298744 9460 298796 9512
rect 356704 9460 356756 9512
rect 471060 9460 471112 9512
rect 291384 9392 291436 9444
rect 421564 9392 421616 9444
rect 190828 9324 190880 9376
rect 283012 9324 283064 9376
rect 368480 9324 368532 9376
rect 524236 9324 524288 9376
rect 222292 9256 222344 9308
rect 402520 9256 402572 9308
rect 222200 9188 222252 9240
rect 406016 9188 406068 9240
rect 223580 9120 223632 9172
rect 409604 9120 409656 9172
rect 79324 9052 79376 9104
rect 90364 9052 90416 9104
rect 95148 9052 95200 9104
rect 107752 9052 107804 9104
rect 226340 9052 226392 9104
rect 420184 9052 420236 9104
rect 56048 8984 56100 9036
rect 98000 8984 98052 9036
rect 164332 8984 164384 9036
rect 179052 8984 179104 9036
rect 227812 8984 227864 9036
rect 423772 8984 423824 9036
rect 424324 8984 424376 9036
rect 480536 8984 480588 9036
rect 482284 8984 482336 9036
rect 497096 8984 497148 9036
rect 12348 8916 12400 8968
rect 57980 8916 58032 8968
rect 71504 8916 71556 8968
rect 130384 8916 130436 8968
rect 173164 8916 173216 8968
rect 203892 8916 203944 8968
rect 230480 8916 230532 8968
rect 437940 8916 437992 8968
rect 483020 8916 483072 8968
rect 514760 8916 514812 8968
rect 428464 8304 428516 8356
rect 434444 8304 434496 8356
rect 74632 8236 74684 8288
rect 83280 8236 83332 8288
rect 224224 8236 224276 8288
rect 225144 8236 225196 8288
rect 258264 8236 258316 8288
rect 300124 8236 300176 8288
rect 332600 8236 332652 8288
rect 382372 8236 382424 8288
rect 244096 8168 244148 8220
rect 296812 8168 296864 8220
rect 333980 8168 334032 8220
rect 385960 8168 386012 8220
rect 282092 8100 282144 8152
rect 422300 8100 422352 8152
rect 242164 8032 242216 8084
rect 303160 8032 303212 8084
rect 375380 8032 375432 8084
rect 549076 8032 549128 8084
rect 199384 7964 199436 8016
rect 274824 7964 274876 8016
rect 376852 7964 376904 8016
rect 552664 7964 552716 8016
rect 205088 7896 205140 7948
rect 287060 7896 287112 7948
rect 328552 7896 328604 7948
rect 368204 7896 368256 7948
rect 376944 7896 376996 7948
rect 556160 7896 556212 7948
rect 187332 7828 187384 7880
rect 282184 7828 282236 7880
rect 329840 7828 329892 7880
rect 371700 7828 371752 7880
rect 378140 7828 378192 7880
rect 559748 7828 559800 7880
rect 176752 7760 176804 7812
rect 280160 7760 280212 7812
rect 297272 7760 297324 7812
rect 310520 7760 310572 7812
rect 331220 7760 331272 7812
rect 375288 7760 375340 7812
rect 380900 7760 380952 7812
rect 570328 7760 570380 7812
rect 80060 7692 80112 7744
rect 104532 7692 104584 7744
rect 200120 7692 200172 7744
rect 320916 7692 320968 7744
rect 331312 7692 331364 7744
rect 378876 7692 378928 7744
rect 382464 7692 382516 7744
rect 573916 7692 573968 7744
rect 26516 7624 26568 7676
rect 60740 7624 60792 7676
rect 62028 7624 62080 7676
rect 70492 7624 70544 7676
rect 78588 7624 78640 7676
rect 132500 7624 132552 7676
rect 136456 7624 136508 7676
rect 153200 7624 153252 7676
rect 162952 7624 163004 7676
rect 175464 7624 175516 7676
rect 175924 7624 175976 7676
rect 189724 7624 189776 7676
rect 191104 7624 191156 7676
rect 207388 7624 207440 7676
rect 209780 7624 209832 7676
rect 356336 7624 356388 7676
rect 382280 7624 382332 7676
rect 577412 7624 577464 7676
rect 38384 7556 38436 7608
rect 93124 7556 93176 7608
rect 114652 7556 114704 7608
rect 123484 7556 123536 7608
rect 131764 7556 131816 7608
rect 385040 7556 385092 7608
rect 356060 7488 356112 7540
rect 387800 7488 387852 7540
rect 279516 6808 279568 6860
rect 306380 6808 306432 6860
rect 318800 6808 318852 6860
rect 329196 6808 329248 6860
rect 337476 6808 337528 6860
rect 403624 6808 403676 6860
rect 305184 6740 305236 6792
rect 386420 6740 386472 6792
rect 266544 6672 266596 6724
rect 367744 6672 367796 6724
rect 187700 6604 187752 6656
rect 267740 6604 267792 6656
rect 276020 6604 276072 6656
rect 305092 6604 305144 6656
rect 320180 6604 320232 6656
rect 332692 6604 332744 6656
rect 357440 6604 357492 6656
rect 481732 6604 481784 6656
rect 187792 6536 187844 6588
rect 271236 6536 271288 6588
rect 272432 6536 272484 6588
rect 305000 6536 305052 6588
rect 320272 6536 320324 6588
rect 336280 6536 336332 6588
rect 358820 6536 358872 6588
rect 485228 6536 485280 6588
rect 190460 6468 190512 6520
rect 281908 6468 281960 6520
rect 321560 6468 321612 6520
rect 339868 6468 339920 6520
rect 360200 6468 360252 6520
rect 488816 6468 488868 6520
rect 191840 6400 191892 6452
rect 285404 6400 285456 6452
rect 286600 6400 286652 6452
rect 307760 6400 307812 6452
rect 322940 6400 322992 6452
rect 343364 6400 343416 6452
rect 363052 6400 363104 6452
rect 499396 6400 499448 6452
rect 191932 6332 191984 6384
rect 288992 6332 289044 6384
rect 290188 6332 290240 6384
rect 309140 6332 309192 6384
rect 323032 6332 323084 6384
rect 346952 6332 347004 6384
rect 362960 6332 363012 6384
rect 502984 6332 503036 6384
rect 91560 6264 91612 6316
rect 106924 6264 106976 6316
rect 193220 6264 193272 6316
rect 292580 6264 292632 6316
rect 293684 6264 293736 6316
rect 309232 6264 309284 6316
rect 324320 6264 324372 6316
rect 350448 6264 350500 6316
rect 364340 6264 364392 6316
rect 506480 6264 506532 6316
rect 81440 6196 81492 6248
rect 108120 6196 108172 6248
rect 129372 6196 129424 6248
rect 151912 6196 151964 6248
rect 194692 6196 194744 6248
rect 296076 6196 296128 6248
rect 327080 6196 327132 6248
rect 361120 6196 361172 6248
rect 365720 6196 365772 6248
rect 510068 6196 510120 6248
rect 512644 6196 512696 6248
rect 525432 6196 525484 6248
rect 572 6128 624 6180
rect 54484 6128 54536 6180
rect 58440 6128 58492 6180
rect 69204 6128 69256 6180
rect 76012 6128 76064 6180
rect 86868 6128 86920 6180
rect 96252 6128 96304 6180
rect 136640 6128 136692 6180
rect 165620 6128 165672 6180
rect 182548 6128 182600 6180
rect 194784 6128 194836 6180
rect 299664 6128 299716 6180
rect 304356 6128 304408 6180
rect 311900 6128 311952 6180
rect 328460 6128 328512 6180
rect 364616 6128 364668 6180
rect 365812 6128 365864 6180
rect 513564 6128 513616 6180
rect 317420 5584 317472 5636
rect 325608 5584 325660 5636
rect 74540 5516 74592 5568
rect 79692 5516 79744 5568
rect 114560 5516 114612 5568
rect 119896 5516 119948 5568
rect 184204 5516 184256 5568
rect 186136 5516 186188 5568
rect 307944 5516 307996 5568
rect 313372 5516 313424 5568
rect 317512 5516 317564 5568
rect 322112 5516 322164 5568
rect 246304 5380 246356 5432
rect 257068 5380 257120 5432
rect 178040 5312 178092 5364
rect 232228 5312 232280 5364
rect 240508 5312 240560 5364
rect 295984 5312 296036 5364
rect 348056 5312 348108 5364
rect 418804 5312 418856 5364
rect 201592 5244 201644 5296
rect 285680 5244 285732 5296
rect 317328 5244 317380 5296
rect 429292 5244 429344 5296
rect 54944 5176 54996 5228
rect 67640 5176 67692 5228
rect 223948 5176 224000 5228
rect 407764 5176 407816 5228
rect 52552 5108 52604 5160
rect 96712 5108 96764 5160
rect 231860 5108 231912 5160
rect 445024 5108 445076 5160
rect 48964 5040 49016 5092
rect 96620 5040 96672 5092
rect 175280 5040 175332 5092
rect 221556 5040 221608 5092
rect 249800 5040 249852 5092
rect 512460 5040 512512 5092
rect 7656 4972 7708 5024
rect 56600 4972 56652 5024
rect 82820 4972 82872 5024
rect 115204 4972 115256 5024
rect 179420 4972 179472 5024
rect 235816 4972 235868 5024
rect 255320 4972 255372 5024
rect 533712 4972 533764 5024
rect 2872 4904 2924 4956
rect 56692 4904 56744 4956
rect 85856 4904 85908 4956
rect 122288 4904 122340 4956
rect 179512 4904 179564 4956
rect 239312 4904 239364 4956
rect 256700 4904 256752 4956
rect 537208 4904 537260 4956
rect 8760 4836 8812 4888
rect 86960 4836 87012 4888
rect 170404 4836 170456 4888
rect 171968 4836 172020 4888
rect 182272 4836 182324 4888
rect 246396 4836 246448 4888
rect 256792 4836 256844 4888
rect 540796 4836 540848 4888
rect 4068 4768 4120 4820
rect 85672 4768 85724 4820
rect 125876 4768 125928 4820
rect 150716 4768 150768 4820
rect 182180 4768 182232 4820
rect 249984 4768 250036 4820
rect 258080 4768 258132 4820
rect 544384 4768 544436 4820
rect 569224 4768 569276 4820
rect 579804 4768 579856 4820
rect 65524 4156 65576 4208
rect 70400 4156 70452 4208
rect 161480 4156 161532 4208
rect 168472 4156 168524 4208
rect 448612 4156 448664 4208
rect 449992 4156 450044 4208
rect 46664 4088 46716 4140
rect 124220 4088 124272 4140
rect 376484 4088 376536 4140
rect 385684 4088 385736 4140
rect 422576 4088 422628 4140
rect 459652 4088 459704 4140
rect 491300 4088 491352 4140
rect 550272 4088 550324 4140
rect 43076 4020 43128 4072
rect 122932 4020 122984 4072
rect 362316 4020 362368 4072
rect 378784 4020 378836 4072
rect 39580 3952 39632 4004
rect 122840 3952 122892 4004
rect 333888 3952 333940 4004
rect 342904 3952 342956 4004
rect 355232 3952 355284 4004
rect 376024 3952 376076 4004
rect 379980 3952 380032 4004
rect 411904 4020 411956 4072
rect 418988 4020 419040 4072
rect 458180 4020 458232 4072
rect 492772 4020 492824 4072
rect 553768 4020 553820 4072
rect 415492 3952 415544 4004
rect 456800 3952 456852 4004
rect 494152 3952 494204 4004
rect 557356 3952 557408 4004
rect 35992 3884 36044 3936
rect 121552 3884 121604 3936
rect 140044 3884 140096 3936
rect 154764 3884 154816 3936
rect 251180 3884 251232 3936
rect 252376 3884 252428 3936
rect 262956 3884 263008 3936
rect 273904 3884 273956 3936
rect 305552 3884 305604 3936
rect 312544 3884 312596 3936
rect 319720 3884 319772 3936
rect 330484 3884 330536 3936
rect 340972 3884 341024 3936
rect 353944 3884 353996 3936
rect 372896 3884 372948 3936
rect 405004 3884 405056 3936
rect 411904 3884 411956 3936
rect 456984 3884 457036 3936
rect 494060 3884 494112 3936
rect 560852 3884 560904 3936
rect 32404 3816 32456 3868
rect 120172 3816 120224 3868
rect 124680 3816 124732 3868
rect 145012 3816 145064 3868
rect 176660 3816 176712 3868
rect 177856 3816 177908 3868
rect 193220 3816 193272 3868
rect 193404 3816 193456 3868
rect 209872 3816 209924 3868
rect 210976 3816 211028 3868
rect 226432 3816 226484 3868
rect 227536 3816 227588 3868
rect 234620 3816 234672 3868
rect 269764 3816 269816 3868
rect 277124 3816 277176 3868
rect 282092 3816 282144 3868
rect 287796 3816 287848 3868
rect 294604 3816 294656 3868
rect 309048 3816 309100 3868
rect 317328 3816 317380 3868
rect 330392 3816 330444 3868
rect 341524 3816 341576 3868
rect 344560 3816 344612 3868
rect 360844 3816 360896 3868
rect 365812 3816 365864 3868
rect 400680 3816 400732 3868
rect 408408 3816 408460 3868
rect 455420 3816 455472 3868
rect 495440 3816 495492 3868
rect 564440 3816 564492 3868
rect 28908 3748 28960 3800
rect 120080 3748 120132 3800
rect 142436 3748 142488 3800
rect 305184 3748 305236 3800
rect 312636 3748 312688 3800
rect 322204 3748 322256 3800
rect 323308 3748 323360 3800
rect 336004 3748 336056 3800
rect 351644 3748 351696 3800
rect 367836 3748 367888 3800
rect 369400 3748 369452 3800
rect 403716 3748 403768 3800
rect 404820 3748 404872 3800
rect 454224 3748 454276 3800
rect 496820 3748 496872 3800
rect 568028 3748 568080 3800
rect 24216 3680 24268 3732
rect 118700 3680 118752 3732
rect 121092 3680 121144 3732
rect 143632 3680 143684 3732
rect 145932 3680 145984 3732
rect 356060 3680 356112 3732
rect 358728 3680 358780 3732
rect 381544 3680 381596 3732
rect 387156 3680 387208 3732
rect 448612 3680 448664 3732
rect 448704 3680 448756 3732
rect 449808 3680 449860 3732
rect 496912 3680 496964 3732
rect 571524 3680 571576 3732
rect 117596 3612 117648 3664
rect 142160 3612 142212 3664
rect 147680 3612 147732 3664
rect 160192 3612 160244 3664
rect 392124 3612 392176 3664
rect 401324 3612 401376 3664
rect 454132 3612 454184 3664
rect 474924 3612 474976 3664
rect 482836 3612 482888 3664
rect 498384 3612 498436 3664
rect 575112 3612 575164 3664
rect 25320 3544 25372 3596
rect 154212 3544 154264 3596
rect 155224 3544 155276 3596
rect 156604 3544 156656 3596
rect 390560 3544 390612 3596
rect 397736 3544 397788 3596
rect 452660 3544 452712 3596
rect 464344 3544 464396 3596
rect 474556 3544 474608 3596
rect 474832 3544 474884 3596
rect 486424 3544 486476 3596
rect 499672 3544 499724 3596
rect 502340 3544 502392 3596
rect 582196 3544 582248 3596
rect 1676 3476 1728 3528
rect 4804 3476 4856 3528
rect 20628 3476 20680 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 15936 3408 15988 3460
rect 146392 3408 146444 3460
rect 11152 3340 11204 3392
rect 15844 3340 15896 3392
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 106924 3340 106976 3392
rect 139400 3340 139452 3392
rect 160100 3476 160152 3528
rect 161296 3476 161348 3528
rect 161388 3476 161440 3528
rect 389180 3476 389232 3528
rect 390652 3476 390704 3528
rect 391848 3476 391900 3528
rect 398840 3476 398892 3528
rect 400128 3476 400180 3528
rect 149520 3408 149572 3460
rect 389272 3408 389324 3460
rect 147772 3340 147824 3392
rect 153016 3340 153068 3392
rect 161388 3340 161440 3392
rect 168380 3340 168432 3392
rect 169576 3340 169628 3392
rect 201500 3340 201552 3392
rect 202696 3340 202748 3392
rect 270040 3340 270092 3392
rect 276664 3340 276716 3392
rect 299572 3340 299624 3392
rect 300768 3340 300820 3392
rect 316132 3340 316184 3392
rect 317328 3340 317380 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 390652 3340 390704 3392
rect 110512 3272 110564 3324
rect 140780 3272 140832 3324
rect 394240 3340 394292 3392
rect 451372 3476 451424 3528
rect 458088 3476 458140 3528
rect 467932 3476 467984 3528
rect 476120 3476 476172 3528
rect 489920 3476 489972 3528
rect 578608 3476 578660 3528
rect 451280 3408 451332 3460
rect 461676 3408 461728 3460
rect 478144 3408 478196 3460
rect 500960 3408 501012 3460
rect 581000 3408 581052 3460
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 426164 3340 426216 3392
rect 459560 3340 459612 3392
rect 491392 3340 491444 3392
rect 546684 3340 546736 3392
rect 433248 3272 433300 3324
rect 462504 3272 462556 3324
rect 490012 3272 490064 3324
rect 543188 3272 543240 3324
rect 13544 3204 13596 3256
rect 14464 3204 14516 3256
rect 114008 3204 114060 3256
rect 142252 3204 142304 3256
rect 440332 3204 440384 3256
rect 441528 3204 441580 3256
rect 443828 3204 443880 3256
rect 465080 3204 465132 3256
rect 488540 3204 488592 3256
rect 539600 3204 539652 3256
rect 19432 3136 19484 3188
rect 117504 3136 117556 3188
rect 280712 3136 280764 3188
rect 284944 3136 284996 3188
rect 531320 3136 531372 3188
rect 532148 3136 532200 3188
rect 316040 3068 316092 3120
rect 318524 3068 318576 3120
rect 316224 3000 316276 3052
rect 324964 3000 325016 3052
rect 473360 3000 473412 3052
rect 479340 3000 479392 3052
rect 9956 2932 10008 2984
rect 11704 2932 11756 2984
rect 298468 2864 298520 2916
rect 304264 2864 304316 2916
rect 199108 2320 199160 2372
rect 401600 2320 401652 2372
rect 192024 2252 192076 2304
rect 400404 2252 400456 2304
rect 181444 2184 181496 2236
rect 396724 2184 396776 2236
rect 167184 2116 167236 2168
rect 393320 2116 393372 2168
rect 237380 2048 237432 2100
rect 466276 2048 466328 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 55445 29866 55473 30048
rect 55324 29838 55473 29866
rect 55836 29866 55864 30049
rect 56600 29912 56652 29918
rect 55836 29838 55904 29866
rect 56754 29866 56782 30049
rect 57655 29918 57683 30049
rect 56600 29854 56652 29860
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 4804 25628 4856 25634
rect 4804 25570 4856 25576
rect 572 6180 624 6186
rect 572 6122 624 6128
rect 584 480 612 6122
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1688 480 1716 3470
rect 2884 480 2912 4898
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 480 4108 4762
rect 4816 3534 4844 25570
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8760 4888 8812 4894
rect 8760 4830 8812 4836
rect 8772 480 8800 4830
rect 10336 3466 10364 26862
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13832 16574 13860 24074
rect 13832 16546 14320 16574
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9968 480 9996 2926
rect 11164 480 11192 3334
rect 11716 2990 11744 15846
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 12360 480 12388 8910
rect 13544 3256 13596 3262
rect 13544 3198 13596 3204
rect 13556 480 13584 3198
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14476 3262 14504 14418
rect 15856 3398 15884 26930
rect 54484 26308 54536 26314
rect 54484 26250 54536 26256
rect 27620 25560 27672 25566
rect 27620 25502 27672 25508
rect 22100 22772 22152 22778
rect 22100 22714 22152 22720
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16592 16574 16620 21422
rect 20720 20188 20772 20194
rect 20720 20130 20772 20136
rect 20732 16574 20760 20130
rect 22112 16574 22140 22714
rect 27632 16574 27660 25502
rect 46940 24268 46992 24274
rect 46940 24210 46992 24216
rect 44180 24200 44232 24206
rect 44180 24142 44232 24148
rect 34520 21412 34572 21418
rect 34520 21354 34572 21360
rect 29000 18896 29052 18902
rect 29000 18838 29052 18844
rect 29012 16574 29040 18838
rect 16592 16546 17080 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 14464 3256 14516 3262
rect 14464 3198 14516 3204
rect 15948 480 15976 3402
rect 17052 480 17080 16546
rect 17960 13116 18012 13122
rect 17960 13058 18012 13064
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 13058
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19444 480 19472 3130
rect 20640 480 20668 3470
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 26516 7676 26568 7682
rect 26516 7618 26568 7624
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24228 480 24256 3674
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 480 25360 3538
rect 26528 480 26556 7618
rect 27724 480 27752 16546
rect 28908 3800 28960 3806
rect 28908 3742 28960 3748
rect 28920 480 28948 3742
rect 30116 480 30144 16546
rect 30840 11756 30892 11762
rect 30840 11698 30892 11704
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 11698
rect 33600 10396 33652 10402
rect 33600 10338 33652 10344
rect 32404 3868 32456 3874
rect 32404 3810 32456 3816
rect 32416 480 32444 3810
rect 33612 480 33640 10338
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 21354
rect 35900 17332 35952 17338
rect 35900 17274 35952 17280
rect 35912 16574 35940 17274
rect 41420 17264 41472 17270
rect 41420 17206 41472 17212
rect 41432 16574 41460 17206
rect 35912 16546 36768 16574
rect 41432 16546 41920 16574
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36004 480 36032 3878
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 40224 15972 40276 15978
rect 40224 15914 40276 15920
rect 38384 7608 38436 7614
rect 38384 7550 38436 7556
rect 38396 480 38424 7550
rect 39580 4004 39632 4010
rect 39580 3946 39632 3952
rect 39592 480 39620 3946
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 15914
rect 41892 480 41920 16546
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43088 480 43116 4014
rect 44192 3398 44220 24142
rect 46952 16574 46980 24210
rect 51080 22976 51132 22982
rect 51080 22918 51132 22924
rect 49700 18624 49752 18630
rect 49700 18566 49752 18572
rect 49712 16574 49740 18566
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44272 11824 44324 11830
rect 44272 11766 44324 11772
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44284 480 44312 11766
rect 46664 4140 46716 4146
rect 46664 4082 46716 4088
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 4082
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 5092 49016 5098
rect 48964 5034 49016 5040
rect 48976 480 49004 5034
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 22918
rect 52460 19984 52512 19990
rect 52460 19926 52512 19932
rect 52472 16574 52500 19926
rect 52472 16546 53328 16574
rect 52552 5160 52604 5166
rect 52552 5102 52604 5108
rect 52564 480 52592 5102
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54496 6186 54524 26250
rect 55324 25634 55352 29838
rect 55876 26314 55904 29838
rect 55864 26308 55916 26314
rect 55864 26250 55916 26256
rect 55312 25628 55364 25634
rect 55312 25570 55364 25576
rect 56048 9036 56100 9042
rect 56048 8978 56100 8984
rect 54484 6180 54536 6186
rect 54484 6122 54536 6128
rect 54944 5228 54996 5234
rect 54944 5170 54996 5176
rect 54956 480 54984 5170
rect 56060 480 56088 8978
rect 56612 5030 56640 29854
rect 56704 29838 56782 29866
rect 57643 29912 57695 29918
rect 58573 29866 58601 30049
rect 59491 29866 59519 30049
rect 60392 29866 60420 30049
rect 61310 29866 61338 30049
rect 57643 29854 57695 29860
rect 57992 29838 58601 29866
rect 59372 29838 59519 29866
rect 60384 29838 60420 29866
rect 61304 29838 61338 29866
rect 62120 29912 62172 29918
rect 62120 29854 62172 29860
rect 62211 29866 62239 30049
rect 63112 29918 63140 30049
rect 63100 29912 63152 29918
rect 56600 5024 56652 5030
rect 56600 4966 56652 4972
rect 56704 4962 56732 29838
rect 56784 10328 56836 10334
rect 56784 10270 56836 10276
rect 56692 4956 56744 4962
rect 56692 4898 56744 4904
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 10270
rect 57992 8974 58020 29838
rect 59372 26234 59400 29838
rect 60384 26234 60412 29838
rect 61304 26234 61332 29838
rect 59280 26206 59400 26234
rect 59464 26206 60412 26234
rect 60752 26206 61332 26234
rect 59280 21486 59308 26206
rect 59268 21480 59320 21486
rect 59268 21422 59320 21428
rect 59464 20194 59492 26206
rect 59452 20188 59504 20194
rect 59452 20130 59504 20136
rect 59360 20052 59412 20058
rect 59360 19994 59412 20000
rect 57980 8968 58032 8974
rect 57980 8910 58032 8916
rect 58440 6180 58492 6186
rect 58440 6122 58492 6128
rect 58452 480 58480 6122
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 19994
rect 60752 7682 60780 26206
rect 60832 14544 60884 14550
rect 60832 14486 60884 14492
rect 60740 7676 60792 7682
rect 60740 7618 60792 7624
rect 60844 480 60872 14486
rect 62132 10402 62160 29854
rect 62211 29838 62252 29866
rect 64013 29866 64041 30049
rect 63100 29854 63152 29860
rect 62224 18902 62252 29838
rect 63512 29838 64041 29866
rect 64931 29866 64959 30049
rect 65815 29866 65843 30049
rect 66750 29866 66778 30049
rect 64931 29838 65012 29866
rect 62212 18896 62264 18902
rect 62212 18838 62264 18844
rect 62212 18760 62264 18766
rect 62212 18702 62264 18708
rect 62224 16574 62252 18702
rect 63512 17338 63540 29838
rect 64880 28144 64932 28150
rect 64880 28086 64932 28092
rect 63500 17332 63552 17338
rect 63500 17274 63552 17280
rect 62224 16546 63264 16574
rect 62120 10396 62172 10402
rect 62120 10338 62172 10344
rect 62028 7676 62080 7682
rect 62028 7618 62080 7624
rect 62040 480 62068 7618
rect 63236 480 63264 16546
rect 64328 13184 64380 13190
rect 64328 13126 64380 13132
rect 64340 480 64368 13126
rect 64892 11830 64920 28086
rect 64984 15978 65012 29838
rect 65812 29838 65843 29866
rect 66732 29838 66778 29866
rect 67634 29866 67662 30049
rect 68569 29866 68597 30049
rect 69453 29866 69481 30049
rect 67634 29838 67772 29866
rect 68569 29838 68600 29866
rect 65812 28150 65840 29838
rect 65800 28144 65852 28150
rect 65800 28086 65852 28092
rect 66732 26234 66760 29838
rect 67640 28144 67692 28150
rect 67640 28086 67692 28092
rect 66272 26206 66760 26234
rect 66272 24274 66300 26206
rect 66260 24268 66312 24274
rect 66260 24210 66312 24216
rect 64972 15972 65024 15978
rect 64972 15914 65024 15920
rect 66720 15972 66772 15978
rect 66720 15914 66772 15920
rect 64880 11824 64932 11830
rect 64880 11766 64932 11772
rect 65524 4208 65576 4214
rect 65524 4150 65576 4156
rect 65536 480 65564 4150
rect 66732 480 66760 15914
rect 67652 5234 67680 28086
rect 67744 22982 67772 29838
rect 68572 28150 68600 29838
rect 69216 29838 69481 29866
rect 68560 28144 68612 28150
rect 68560 28086 68612 28092
rect 69020 27600 69072 27606
rect 69020 27542 69072 27548
rect 67732 22976 67784 22982
rect 67732 22918 67784 22924
rect 67732 22840 67784 22846
rect 67732 22782 67784 22788
rect 67640 5228 67692 5234
rect 67640 5170 67692 5176
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67744 354 67772 22782
rect 69032 3482 69060 27542
rect 69112 24268 69164 24274
rect 69112 24210 69164 24216
rect 69124 3618 69152 24210
rect 69216 6186 69244 29838
rect 70388 29832 70416 30049
rect 71289 29832 71317 30049
rect 70388 29804 70532 29832
rect 70400 26104 70452 26110
rect 70400 26046 70452 26052
rect 69204 6180 69256 6186
rect 69204 6122 69256 6128
rect 70412 4214 70440 26046
rect 70504 7682 70532 29804
rect 71240 29804 71317 29832
rect 71872 29844 71924 29850
rect 71240 26110 71268 29804
rect 72207 29832 72235 30049
rect 73091 29850 73119 30049
rect 74043 29866 74071 30049
rect 71872 29786 71924 29792
rect 72160 29804 72235 29832
rect 73079 29844 73131 29850
rect 71228 26104 71280 26110
rect 71228 26046 71280 26052
rect 71884 16574 71912 29786
rect 72160 27606 72188 29804
rect 74043 29838 74120 29866
rect 73079 29786 73131 29792
rect 72148 27600 72200 27606
rect 72148 27542 72200 27548
rect 74092 26314 74120 29838
rect 74910 29832 74938 30049
rect 75845 29832 75873 30049
rect 76746 29832 76774 30049
rect 74552 29804 74938 29832
rect 75840 29804 75873 29832
rect 76668 29804 76774 29832
rect 77300 29844 77352 29850
rect 74080 26308 74132 26314
rect 74080 26250 74132 26256
rect 73160 17400 73212 17406
rect 73160 17342 73212 17348
rect 73172 16574 73200 17342
rect 71884 16546 72648 16574
rect 73172 16546 73384 16574
rect 71504 8968 71556 8974
rect 71504 8910 71556 8916
rect 70492 7676 70544 7682
rect 70492 7618 70544 7624
rect 70400 4208 70452 4214
rect 70400 4150 70452 4156
rect 69124 3590 69888 3618
rect 69032 3454 69152 3482
rect 69124 480 69152 3454
rect 67886 354 67998 480
rect 67744 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 3590
rect 71516 480 71544 8910
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 74552 5574 74580 29804
rect 75840 26110 75868 29804
rect 75920 26308 75972 26314
rect 75920 26250 75972 26256
rect 74632 26104 74684 26110
rect 74632 26046 74684 26052
rect 75828 26104 75880 26110
rect 75828 26046 75880 26052
rect 74644 8294 74672 26046
rect 74724 21480 74776 21486
rect 74724 21422 74776 21428
rect 74736 16574 74764 21422
rect 74736 16546 75040 16574
rect 74632 8288 74684 8294
rect 74632 8230 74684 8236
rect 74540 5568 74592 5574
rect 74540 5510 74592 5516
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 26250
rect 76668 22094 76696 29804
rect 77647 29832 77675 30049
rect 78565 29850 78593 30049
rect 78553 29844 78605 29850
rect 77647 29804 77708 29832
rect 77300 29786 77352 29792
rect 76024 22066 76696 22094
rect 76024 6186 76052 22066
rect 77312 11966 77340 29786
rect 77680 26382 77708 29804
rect 79466 29832 79494 30049
rect 80384 29866 80412 30049
rect 78553 29786 78605 29792
rect 79428 29804 79494 29832
rect 80060 29844 80112 29850
rect 79428 26874 79456 29804
rect 80060 29786 80112 29792
rect 80348 29838 80412 29866
rect 81302 29850 81330 30049
rect 82203 29866 82231 30049
rect 83121 29866 83149 30049
rect 81290 29844 81342 29850
rect 79244 26846 79456 26874
rect 77668 26376 77720 26382
rect 77668 26318 77720 26324
rect 79244 22094 79272 26846
rect 79324 26376 79376 26382
rect 79324 26318 79376 26324
rect 78692 22066 79272 22094
rect 77300 11960 77352 11966
rect 77300 11902 77352 11908
rect 77392 10464 77444 10470
rect 77392 10406 77444 10412
rect 76012 6180 76064 6186
rect 76012 6122 76064 6128
rect 77404 480 77432 10406
rect 78692 10402 78720 22066
rect 78680 10396 78732 10402
rect 78680 10338 78732 10344
rect 79336 9110 79364 26318
rect 79324 9104 79376 9110
rect 79324 9046 79376 9052
rect 80072 7750 80100 29786
rect 80348 26234 80376 29838
rect 81290 29786 81342 29792
rect 81452 29838 82231 29866
rect 82820 29844 82872 29850
rect 80256 26206 80376 26234
rect 80152 21548 80204 21554
rect 80152 21490 80204 21496
rect 80060 7744 80112 7750
rect 80060 7686 80112 7692
rect 78588 7676 78640 7682
rect 78588 7618 78640 7624
rect 78600 480 78628 7618
rect 80164 6914 80192 21490
rect 80256 13258 80284 26206
rect 80244 13252 80296 13258
rect 80244 13194 80296 13200
rect 80164 6886 80928 6914
rect 79692 5568 79744 5574
rect 79692 5510 79744 5516
rect 79704 480 79732 5510
rect 80900 480 80928 6886
rect 81452 6254 81480 29838
rect 82820 29786 82872 29792
rect 82924 29838 83149 29866
rect 84005 29850 84033 30049
rect 83993 29844 84045 29850
rect 81532 17332 81584 17338
rect 81532 17274 81584 17280
rect 81544 16574 81572 17274
rect 81544 16546 81664 16574
rect 81440 6248 81492 6254
rect 81440 6190 81492 6196
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 82832 5030 82860 29786
rect 82924 14618 82952 29838
rect 84923 29832 84951 30049
rect 83993 29786 84045 29792
rect 84212 29804 84951 29832
rect 85672 29844 85724 29850
rect 84212 25702 84240 29804
rect 85841 29832 85869 30049
rect 86742 29850 86770 30049
rect 86730 29844 86782 29850
rect 85841 29804 85896 29832
rect 85672 29786 85724 29792
rect 84200 25696 84252 25702
rect 84200 25638 84252 25644
rect 82912 14612 82964 14618
rect 82912 14554 82964 14560
rect 84200 11892 84252 11898
rect 84200 11834 84252 11840
rect 83280 8288 83332 8294
rect 83280 8230 83332 8236
rect 82820 5024 82872 5030
rect 82820 4966 82872 4972
rect 83292 480 83320 8230
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 11834
rect 85684 4826 85712 29786
rect 85764 11824 85816 11830
rect 85764 11766 85816 11772
rect 85672 4820 85724 4826
rect 85672 4762 85724 4768
rect 85776 3482 85804 11766
rect 85868 4962 85896 29804
rect 87660 29832 87688 30049
rect 86730 29786 86782 29792
rect 87616 29804 87688 29832
rect 88432 29844 88484 29850
rect 87616 26234 87644 29804
rect 88578 29832 88606 30049
rect 89462 29850 89490 30049
rect 88432 29786 88484 29792
rect 88536 29804 88606 29832
rect 89450 29844 89502 29850
rect 86972 26206 87644 26234
rect 86868 6180 86920 6186
rect 86868 6122 86920 6128
rect 85856 4956 85908 4962
rect 85856 4898 85908 4904
rect 85684 3454 85804 3482
rect 85684 480 85712 3454
rect 86880 480 86908 6122
rect 86972 4894 87000 26206
rect 88340 25628 88392 25634
rect 88340 25570 88392 25576
rect 87052 22908 87104 22914
rect 87052 22850 87104 22856
rect 87064 16574 87092 22850
rect 87064 16546 87552 16574
rect 86960 4888 87012 4894
rect 86960 4830 87012 4836
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 88352 6914 88380 25570
rect 88444 13122 88472 29786
rect 88536 14482 88564 29804
rect 90397 29832 90425 30049
rect 91281 29832 91309 30049
rect 89450 29786 89502 29792
rect 89732 29804 90425 29832
rect 91204 29804 91309 29832
rect 89732 22778 89760 29804
rect 90364 27600 90416 27606
rect 90364 27542 90416 27548
rect 89720 22772 89772 22778
rect 89720 22714 89772 22720
rect 88524 14476 88576 14482
rect 88524 14418 88576 14424
rect 88432 13116 88484 13122
rect 88432 13058 88484 13064
rect 90376 11762 90404 27542
rect 91204 26234 91232 29804
rect 92216 27606 92244 30049
rect 93117 29832 93145 30049
rect 94035 29866 94063 30049
rect 94936 29866 94964 30049
rect 95837 29866 95865 30049
rect 96738 29866 96766 30049
rect 97673 29866 97701 30049
rect 98557 29866 98585 30049
rect 99492 29866 99520 30049
rect 100393 29866 100421 30049
rect 101294 29866 101322 30049
rect 94035 29838 94084 29866
rect 92492 29804 93145 29832
rect 92204 27600 92256 27606
rect 92204 27542 92256 27548
rect 91020 26206 91232 26234
rect 91020 25566 91048 26206
rect 91008 25560 91060 25566
rect 91008 25502 91060 25508
rect 92492 21418 92520 29804
rect 94056 26382 94084 29838
rect 94884 29838 94964 29866
rect 95804 29838 95865 29866
rect 96632 29838 96766 29866
rect 96816 29838 97701 29866
rect 98012 29838 98585 29866
rect 99392 29838 99520 29866
rect 99852 29838 100421 29866
rect 101232 29838 101322 29866
rect 102212 29866 102240 30049
rect 103113 29866 103141 30049
rect 104031 29866 104059 30049
rect 102212 29838 102272 29866
rect 93124 26376 93176 26382
rect 93124 26318 93176 26324
rect 94044 26376 94096 26382
rect 94044 26318 94096 26324
rect 92480 21412 92532 21418
rect 92480 21354 92532 21360
rect 92480 18692 92532 18698
rect 92480 18634 92532 18640
rect 90364 11756 90416 11762
rect 90364 11698 90416 11704
rect 90364 9104 90416 9110
rect 90364 9046 90416 9052
rect 88352 6886 89208 6914
rect 89180 480 89208 6886
rect 90376 480 90404 9046
rect 91560 6316 91612 6322
rect 91560 6258 91612 6264
rect 91572 480 91600 6258
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 18634
rect 93136 7614 93164 26318
rect 94884 26234 94912 29838
rect 95804 27266 95832 29838
rect 95148 27260 95200 27266
rect 95148 27202 95200 27208
rect 95792 27260 95844 27266
rect 95792 27202 95844 27208
rect 93964 26206 94912 26234
rect 93964 17270 93992 26206
rect 95160 24206 95188 27202
rect 95148 24200 95200 24206
rect 95148 24142 95200 24148
rect 93952 17264 94004 17270
rect 93952 17206 94004 17212
rect 93952 11960 94004 11966
rect 93952 11902 94004 11908
rect 93124 7608 93176 7614
rect 93124 7550 93176 7556
rect 93964 480 93992 11902
rect 95148 9104 95200 9110
rect 95148 9046 95200 9052
rect 95160 480 95188 9046
rect 96252 6180 96304 6186
rect 96252 6122 96304 6128
rect 96264 480 96292 6122
rect 96632 5098 96660 29838
rect 96816 26234 96844 29838
rect 96724 26206 96844 26234
rect 96724 5166 96752 26206
rect 97448 10396 97500 10402
rect 97448 10338 97500 10344
rect 96712 5160 96764 5166
rect 96712 5102 96764 5108
rect 96620 5092 96672 5098
rect 96620 5034 96672 5040
rect 97460 480 97488 10338
rect 98012 9042 98040 29838
rect 99392 26234 99420 29838
rect 99852 26234 99880 29838
rect 101232 26234 101260 29838
rect 102140 28144 102192 28150
rect 102140 28086 102192 28092
rect 99300 26206 99420 26234
rect 99484 26206 99880 26234
rect 100772 26206 101260 26234
rect 98092 20120 98144 20126
rect 98092 20062 98144 20068
rect 98104 16574 98132 20062
rect 99300 20058 99328 26206
rect 99380 24200 99432 24206
rect 99380 24142 99432 24148
rect 99288 20052 99340 20058
rect 99288 19994 99340 20000
rect 99392 16574 99420 24142
rect 99484 18766 99512 26206
rect 99472 18760 99524 18766
rect 99472 18702 99524 18708
rect 98104 16546 98224 16574
rect 99392 16546 99880 16574
rect 98000 9036 98052 9042
rect 98000 8978 98052 8984
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 100772 15978 100800 26206
rect 102152 17406 102180 28086
rect 102244 24274 102272 29838
rect 103072 29838 103141 29866
rect 103532 29838 104059 29866
rect 104949 29866 104977 30049
rect 105850 29866 105878 30049
rect 106768 29866 106796 30049
rect 104949 29838 105032 29866
rect 103072 28150 103100 29838
rect 103060 28144 103112 28150
rect 103060 28086 103112 28092
rect 102232 24268 102284 24274
rect 102232 24210 102284 24216
rect 102140 17400 102192 17406
rect 102140 17342 102192 17348
rect 100760 15972 100812 15978
rect 100760 15914 100812 15920
rect 102232 15972 102284 15978
rect 102232 15914 102284 15920
rect 100760 13252 100812 13258
rect 100760 13194 100812 13200
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 13194
rect 102244 480 102272 15914
rect 103532 10470 103560 29838
rect 104900 28144 104952 28150
rect 104900 28086 104952 28092
rect 104912 11898 104940 28086
rect 105004 21554 105032 29838
rect 105832 29838 105878 29866
rect 106752 29838 106796 29866
rect 107652 29866 107680 30049
rect 108570 29866 108598 30049
rect 107652 29838 107700 29866
rect 105832 28150 105860 29838
rect 105820 28144 105872 28150
rect 105820 28086 105872 28092
rect 106752 26234 106780 29838
rect 107672 27606 107700 29838
rect 108500 29838 108598 29866
rect 109488 29866 109516 30049
rect 110389 29866 110417 30049
rect 111307 29866 111335 30049
rect 112225 29866 112253 30049
rect 109488 29838 109540 29866
rect 110389 29838 110552 29866
rect 106924 27600 106976 27606
rect 106924 27542 106976 27548
rect 107660 27600 107712 27606
rect 107660 27542 107712 27548
rect 106292 26206 106780 26234
rect 106292 22914 106320 26206
rect 106280 22908 106332 22914
rect 106280 22850 106332 22856
rect 104992 21548 105044 21554
rect 104992 21490 105044 21496
rect 105728 12504 105780 12510
rect 105728 12446 105780 12452
rect 104900 11892 104952 11898
rect 104900 11834 104952 11840
rect 103520 10464 103572 10470
rect 103520 10406 103572 10412
rect 103336 10396 103388 10402
rect 103336 10338 103388 10344
rect 103348 480 103376 10338
rect 104532 7744 104584 7750
rect 104532 7686 104584 7692
rect 104544 480 104572 7686
rect 105740 480 105768 12446
rect 106936 6322 106964 27542
rect 108500 26234 108528 29838
rect 109512 27606 109540 29838
rect 110420 28144 110472 28150
rect 110420 28086 110472 28092
rect 108948 27600 109000 27606
rect 108948 27542 109000 27548
rect 109500 27600 109552 27606
rect 109500 27542 109552 27548
rect 107764 26206 108528 26234
rect 107764 9110 107792 26206
rect 108960 20126 108988 27542
rect 109040 27532 109092 27538
rect 109040 27474 109092 27480
rect 108948 20120 109000 20126
rect 108948 20062 109000 20068
rect 107752 9104 107804 9110
rect 107752 9046 107804 9052
rect 106924 6316 106976 6322
rect 106924 6258 106976 6264
rect 108120 6248 108172 6254
rect 108120 6190 108172 6196
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 106936 480 106964 3334
rect 108132 480 108160 6190
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 27474
rect 110432 12510 110460 28086
rect 110524 15978 110552 29838
rect 111260 29838 111335 29866
rect 111892 29844 111944 29850
rect 111260 28150 111288 29838
rect 111892 29786 111944 29792
rect 112180 29838 112253 29866
rect 113109 29850 113137 30049
rect 114044 29866 114072 30049
rect 114928 29866 114956 30049
rect 115863 29866 115891 30049
rect 116764 29866 116792 30049
rect 113097 29844 113149 29850
rect 111248 28144 111300 28150
rect 111248 28086 111300 28092
rect 111904 16574 111932 29786
rect 112180 27538 112208 29838
rect 113097 29786 113149 29792
rect 114020 29838 114072 29866
rect 114572 29838 114956 29866
rect 115860 29838 115891 29866
rect 116688 29838 116792 29866
rect 117682 29866 117710 30049
rect 118566 29866 118594 30049
rect 119518 29866 119546 30049
rect 120385 29866 120413 30049
rect 121320 29866 121348 30049
rect 122204 29866 122232 30049
rect 123139 29866 123167 30049
rect 124040 29866 124068 30049
rect 124941 29866 124969 30049
rect 125859 29866 125887 30049
rect 126777 29866 126805 30049
rect 127678 29866 127706 30049
rect 128596 29866 128624 30049
rect 117682 29838 117728 29866
rect 114020 27606 114048 29838
rect 114008 27600 114060 27606
rect 114008 27542 114060 27548
rect 112168 27532 112220 27538
rect 112168 27474 112220 27480
rect 111904 16546 112392 16574
rect 110512 15972 110564 15978
rect 110512 15914 110564 15920
rect 111616 14612 111668 14618
rect 111616 14554 111668 14560
rect 110420 12504 110472 12510
rect 110420 12446 110472 12452
rect 110512 3324 110564 3330
rect 110512 3266 110564 3272
rect 110524 480 110552 3266
rect 111628 480 111656 14554
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114572 5574 114600 29838
rect 115860 28150 115888 29838
rect 114652 28144 114704 28150
rect 114652 28086 114704 28092
rect 115848 28144 115900 28150
rect 115848 28086 115900 28092
rect 114664 7614 114692 28086
rect 115940 27600 115992 27606
rect 115940 27542 115992 27548
rect 114652 7608 114704 7614
rect 114652 7550 114704 7556
rect 115952 6914 115980 27542
rect 116688 26234 116716 29838
rect 117700 27606 117728 29838
rect 118528 29838 118594 29866
rect 119448 29838 119546 29866
rect 120092 29838 120413 29866
rect 121288 29838 121348 29866
rect 122116 29838 122232 29866
rect 122852 29838 123167 29866
rect 123956 29838 124068 29866
rect 124232 29838 124969 29866
rect 125612 29838 125887 29866
rect 125980 29838 126805 29866
rect 127636 29838 127706 29866
rect 128360 29844 128412 29850
rect 117228 27600 117280 27606
rect 117228 27542 117280 27548
rect 117688 27600 117740 27606
rect 117688 27542 117740 27548
rect 116044 26206 116716 26234
rect 116044 15910 116072 26206
rect 117240 24138 117268 27542
rect 118528 26234 118556 29838
rect 119448 26234 119476 29838
rect 117516 26206 118556 26234
rect 118712 26206 119476 26234
rect 117228 24132 117280 24138
rect 117228 24074 117280 24080
rect 116032 15904 116084 15910
rect 116032 15846 116084 15852
rect 115952 6886 116440 6914
rect 114560 5568 114612 5574
rect 114560 5510 114612 5516
rect 115204 5024 115256 5030
rect 115204 4966 115256 4972
rect 114008 3256 114060 3262
rect 114008 3198 114060 3204
rect 114020 480 114048 3198
rect 115216 480 115244 4966
rect 116412 480 116440 6886
rect 117516 3194 117544 26206
rect 118712 3738 118740 26206
rect 118792 25696 118844 25702
rect 118792 25638 118844 25644
rect 118700 3732 118752 3738
rect 118700 3674 118752 3680
rect 117596 3664 117648 3670
rect 117596 3606 117648 3612
rect 117504 3188 117556 3194
rect 117504 3130 117556 3136
rect 117608 480 117636 3606
rect 118804 480 118832 25638
rect 119896 5568 119948 5574
rect 119896 5510 119948 5516
rect 119908 480 119936 5510
rect 120092 3806 120120 29838
rect 121288 26234 121316 29838
rect 122116 26234 122144 29838
rect 120184 26206 121316 26234
rect 121564 26206 122144 26234
rect 120184 3874 120212 26206
rect 121564 3942 121592 26206
rect 122288 4956 122340 4962
rect 122288 4898 122340 4904
rect 121552 3936 121604 3942
rect 121552 3878 121604 3884
rect 120172 3868 120224 3874
rect 120172 3810 120224 3816
rect 120080 3800 120132 3806
rect 120080 3742 120132 3748
rect 121092 3732 121144 3738
rect 121092 3674 121144 3680
rect 121104 480 121132 3674
rect 122300 480 122328 4898
rect 122852 4010 122880 29838
rect 123956 26234 123984 29838
rect 122944 26206 123984 26234
rect 122944 4078 122972 26206
rect 123484 7608 123536 7614
rect 123484 7550 123536 7556
rect 122932 4072 122984 4078
rect 122932 4014 122984 4020
rect 122840 4004 122892 4010
rect 122840 3946 122892 3952
rect 123496 480 123524 7550
rect 124232 4146 124260 29838
rect 125612 18630 125640 29838
rect 125980 26234 126008 29838
rect 127636 27606 127664 29838
rect 128360 29786 128412 29792
rect 128556 29838 128624 29866
rect 129497 29850 129525 30049
rect 130398 29866 130426 30049
rect 129485 29844 129537 29850
rect 126244 27600 126296 27606
rect 126244 27542 126296 27548
rect 127624 27600 127676 27606
rect 127624 27542 127676 27548
rect 125704 26206 126008 26234
rect 125704 19990 125732 26206
rect 125692 19984 125744 19990
rect 125692 19926 125744 19932
rect 125600 18624 125652 18630
rect 125600 18566 125652 18572
rect 126256 10334 126284 27542
rect 126980 16108 127032 16114
rect 126980 16050 127032 16056
rect 126244 10328 126296 10334
rect 126244 10270 126296 10276
rect 125876 4820 125928 4826
rect 125876 4762 125928 4768
rect 124220 4140 124272 4146
rect 124220 4082 124272 4088
rect 124680 3868 124732 3874
rect 124680 3810 124732 3816
rect 124692 480 124720 3810
rect 125888 480 125916 4762
rect 126992 480 127020 16050
rect 128372 13190 128400 29786
rect 128556 26234 128584 29838
rect 129485 29786 129537 29792
rect 130304 29838 130426 29866
rect 130304 26234 130332 29838
rect 131333 29730 131361 30049
rect 132217 29866 132245 30049
rect 133135 29866 133163 30049
rect 134036 29866 134064 30049
rect 131316 29702 131361 29730
rect 131408 29838 132245 29866
rect 132512 29838 133163 29866
rect 133880 29844 133932 29850
rect 131316 27198 131344 29702
rect 130384 27192 130436 27198
rect 130384 27134 130436 27140
rect 131304 27192 131356 27198
rect 131304 27134 131356 27140
rect 128464 26206 128584 26234
rect 129752 26206 130332 26234
rect 128464 14550 128492 26206
rect 129752 22846 129780 26206
rect 129832 23044 129884 23050
rect 129832 22986 129884 22992
rect 129740 22840 129792 22846
rect 129740 22782 129792 22788
rect 128452 14544 128504 14550
rect 128452 14486 128504 14492
rect 128360 13184 128412 13190
rect 128360 13126 128412 13132
rect 128176 13116 128228 13122
rect 128176 13058 128228 13064
rect 128188 480 128216 13058
rect 129844 6914 129872 22986
rect 130396 8974 130424 27134
rect 131408 26234 131436 29838
rect 131224 26206 131436 26234
rect 131224 21486 131252 26206
rect 131212 21480 131264 21486
rect 131212 21422 131264 21428
rect 130384 8968 130436 8974
rect 130384 8910 130436 8916
rect 132512 7682 132540 29838
rect 133880 29786 133932 29792
rect 133984 29838 134064 29866
rect 134954 29850 134982 30049
rect 135872 29866 135900 30049
rect 136756 29866 136784 30049
rect 134942 29844 134994 29850
rect 132960 15972 133012 15978
rect 132960 15914 133012 15920
rect 132500 7676 132552 7682
rect 132500 7618 132552 7624
rect 131764 7608 131816 7614
rect 131764 7550 131816 7556
rect 129844 6886 130608 6914
rect 129372 6248 129424 6254
rect 129372 6190 129424 6196
rect 129384 480 129412 6190
rect 130580 480 130608 6886
rect 131776 480 131804 7550
rect 132972 480 133000 15914
rect 133892 11830 133920 29786
rect 133984 17338 134012 29838
rect 134942 29786 134994 29792
rect 135824 29838 135900 29866
rect 136640 29844 136692 29850
rect 135824 26234 135852 29838
rect 136640 29786 136692 29792
rect 136744 29838 136784 29866
rect 137691 29850 137719 30049
rect 138592 29866 138620 30049
rect 139510 29866 139538 30049
rect 137679 29844 137731 29850
rect 135272 26206 135852 26234
rect 135272 25634 135300 26206
rect 135260 25628 135312 25634
rect 135260 25570 135312 25576
rect 133972 17332 134024 17338
rect 133972 17274 134024 17280
rect 135260 14476 135312 14482
rect 135260 14418 135312 14424
rect 133880 11824 133932 11830
rect 133880 11766 133932 11772
rect 133972 11824 134024 11830
rect 133972 11766 134024 11772
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133984 354 134012 11766
rect 135272 480 135300 14418
rect 136456 7676 136508 7682
rect 136456 7618 136508 7624
rect 136468 480 136496 7618
rect 136652 6186 136680 29786
rect 136744 18698 136772 29838
rect 137679 29786 137731 29792
rect 138584 29838 138620 29866
rect 139400 29844 139452 29850
rect 138584 26234 138612 29838
rect 139400 29786 139452 29792
rect 139504 29838 139538 29866
rect 140411 29850 140439 30049
rect 141329 29866 141357 30049
rect 140399 29844 140451 29850
rect 138032 26206 138612 26234
rect 138032 24206 138060 26206
rect 138020 24200 138072 24206
rect 138020 24142 138072 24148
rect 136824 20392 136876 20398
rect 136824 20334 136876 20340
rect 136732 18692 136784 18698
rect 136732 18634 136784 18640
rect 136836 16574 136864 20334
rect 136836 16546 137232 16574
rect 136640 6180 136692 6186
rect 136640 6122 136692 6128
rect 134126 354 134238 480
rect 133984 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138848 15904 138900 15910
rect 138848 15846 138900 15852
rect 138860 480 138888 15846
rect 139412 3398 139440 29786
rect 139504 10402 139532 29838
rect 140399 29786 140451 29792
rect 140792 29838 141357 29866
rect 142213 29866 142241 30049
rect 143165 29866 143193 30049
rect 144032 29866 144060 30049
rect 142213 29838 142292 29866
rect 139492 10396 139544 10402
rect 139492 10338 139544 10344
rect 140044 3936 140096 3942
rect 140044 3878 140096 3884
rect 139400 3392 139452 3398
rect 139400 3334 139452 3340
rect 140056 480 140084 3878
rect 140792 3330 140820 29838
rect 142160 28144 142212 28150
rect 142160 28086 142212 28092
rect 140872 19100 140924 19106
rect 140872 19042 140924 19048
rect 140884 16574 140912 19042
rect 140884 16546 141280 16574
rect 140780 3324 140832 3330
rect 140780 3266 140832 3272
rect 141252 480 141280 16546
rect 142172 3670 142200 28086
rect 142160 3664 142212 3670
rect 142160 3606 142212 3612
rect 142264 3262 142292 29838
rect 143092 29838 143193 29866
rect 144012 29838 144060 29866
rect 144967 29866 144995 30049
rect 145868 29866 145896 30049
rect 146786 29866 146814 30049
rect 144967 29838 145052 29866
rect 143092 28150 143120 29838
rect 143080 28144 143132 28150
rect 143080 28086 143132 28092
rect 143540 27056 143592 27062
rect 143540 26998 143592 27004
rect 142436 3800 142488 3806
rect 142436 3742 142488 3748
rect 142252 3256 142304 3262
rect 142252 3198 142304 3204
rect 142448 480 142476 3742
rect 143552 480 143580 26998
rect 144012 26234 144040 29838
rect 143644 26206 144040 26234
rect 143644 3738 143672 26206
rect 143724 21888 143776 21894
rect 143724 21830 143776 21836
rect 143736 16574 143764 21830
rect 143736 16546 144776 16574
rect 143632 3732 143684 3738
rect 143632 3674 143684 3680
rect 144748 480 144776 16546
rect 145024 3874 145052 29838
rect 145852 29838 145896 29866
rect 146772 29838 146814 29866
rect 147687 29866 147715 30049
rect 148588 29866 148616 30049
rect 147687 29838 147812 29866
rect 145852 26994 145880 29838
rect 145840 26988 145892 26994
rect 145840 26930 145892 26936
rect 146300 26988 146352 26994
rect 146300 26930 146352 26936
rect 145012 3868 145064 3874
rect 145012 3810 145064 3816
rect 145932 3732 145984 3738
rect 145932 3674 145984 3680
rect 145944 480 145972 3674
rect 146312 2774 146340 26930
rect 146772 26234 146800 29838
rect 147680 28144 147732 28150
rect 147680 28086 147732 28092
rect 146404 26206 146800 26234
rect 146404 3466 146432 26206
rect 147692 3670 147720 28086
rect 147680 3664 147732 3670
rect 147680 3606 147732 3612
rect 146392 3460 146444 3466
rect 146392 3402 146444 3408
rect 147784 3398 147812 29838
rect 148520 29838 148616 29866
rect 149506 29866 149534 30049
rect 150424 29866 150452 30049
rect 151325 29866 151353 30049
rect 152243 29866 152271 30049
rect 153127 29866 153155 30049
rect 154045 29866 154073 30049
rect 154963 29866 154991 30049
rect 149506 29838 149560 29866
rect 150424 29838 150572 29866
rect 148520 28150 148548 29838
rect 148508 28144 148560 28150
rect 148508 28086 148560 28092
rect 149532 26926 149560 29838
rect 149520 26920 149572 26926
rect 149520 26862 149572 26868
rect 150440 26920 150492 26926
rect 150440 26862 150492 26868
rect 147864 23180 147916 23186
rect 147864 23122 147916 23128
rect 147772 3392 147824 3398
rect 147772 3334 147824 3340
rect 146312 2746 147168 2774
rect 147140 480 147168 2746
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 23122
rect 150452 3482 150480 26862
rect 150544 3641 150572 29838
rect 150636 29838 151353 29866
rect 151832 29838 152271 29866
rect 153120 29838 153155 29866
rect 153212 29838 154073 29866
rect 154776 29838 154991 29866
rect 155864 29866 155892 30049
rect 156782 29866 156810 30049
rect 157700 29866 157728 30049
rect 158601 29866 158629 30049
rect 159519 29866 159547 30049
rect 160403 29866 160431 30049
rect 161338 29866 161366 30049
rect 162239 29866 162267 30049
rect 163157 29866 163185 30049
rect 164058 29866 164086 30049
rect 164993 29866 165021 30049
rect 165860 29866 165888 30049
rect 155864 29838 155908 29866
rect 156782 29838 156828 29866
rect 157700 29838 157748 29866
rect 150636 16574 150664 29838
rect 150636 16546 150756 16574
rect 150728 4826 150756 16546
rect 151832 6914 151860 29838
rect 153120 28150 153148 29838
rect 151912 28144 151964 28150
rect 151912 28086 151964 28092
rect 153108 28144 153160 28150
rect 153108 28086 153160 28092
rect 151924 15978 151952 28086
rect 151912 15972 151964 15978
rect 151912 15914 151964 15920
rect 152004 13456 152056 13462
rect 152004 13398 152056 13404
rect 151832 6886 151952 6914
rect 151924 6254 151952 6886
rect 151912 6248 151964 6254
rect 151912 6190 151964 6196
rect 150716 4820 150768 4826
rect 150716 4762 150768 4768
rect 150530 3632 150586 3641
rect 150530 3567 150586 3576
rect 152016 3482 152044 13398
rect 153212 7682 153240 29838
rect 154672 13524 154724 13530
rect 154672 13466 154724 13472
rect 153200 7676 153252 7682
rect 153200 7618 153252 7624
rect 154212 3596 154264 3602
rect 154212 3538 154264 3544
rect 149520 3460 149572 3466
rect 150452 3454 150664 3482
rect 149520 3402 149572 3408
rect 149532 480 149560 3402
rect 150636 480 150664 3454
rect 151832 3454 152044 3482
rect 151832 480 151860 3454
rect 153016 3392 153068 3398
rect 153016 3334 153068 3340
rect 153028 480 153056 3334
rect 154224 480 154252 3538
rect 154684 3482 154712 13466
rect 154776 3942 154804 29838
rect 155224 27600 155276 27606
rect 155224 27542 155276 27548
rect 154764 3936 154816 3942
rect 154764 3878 154816 3884
rect 155236 3602 155264 27542
rect 155880 27062 155908 29838
rect 155868 27056 155920 27062
rect 155868 26998 155920 27004
rect 156800 26994 156828 29838
rect 156788 26988 156840 26994
rect 156788 26930 156840 26936
rect 157720 26926 157748 29838
rect 158548 29838 158629 29866
rect 159468 29838 159547 29866
rect 160112 29838 160431 29866
rect 161308 29838 161366 29866
rect 161492 29838 162267 29866
rect 163148 29838 163185 29866
rect 163976 29838 164086 29866
rect 164344 29838 165021 29866
rect 165816 29838 165888 29866
rect 166795 29866 166823 30049
rect 167679 29866 167707 30049
rect 168614 29866 168642 30049
rect 169515 29866 169543 30049
rect 170433 29866 170461 30049
rect 166795 29838 166856 29866
rect 158548 27606 158576 29838
rect 158536 27600 158588 27606
rect 158536 27542 158588 27548
rect 157708 26920 157760 26926
rect 157708 26862 157760 26868
rect 159468 26722 159496 29838
rect 157524 26716 157576 26722
rect 157524 26658 157576 26664
rect 159456 26716 159508 26722
rect 159456 26658 159508 26664
rect 157536 16574 157564 26658
rect 157536 16546 157840 16574
rect 155224 3596 155276 3602
rect 155224 3538 155276 3544
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 154684 3454 155448 3482
rect 155420 480 155448 3454
rect 156616 480 156644 3538
rect 157812 480 157840 16546
rect 158904 13592 158956 13598
rect 158904 13534 158956 13540
rect 158916 480 158944 13534
rect 160112 3534 160140 29838
rect 161308 26926 161336 29838
rect 161296 26920 161348 26926
rect 161296 26862 161348 26868
rect 161492 4214 161520 29838
rect 162860 28280 162912 28286
rect 162860 28222 162912 28228
rect 162032 10464 162084 10470
rect 162032 10406 162084 10412
rect 161480 4208 161532 4214
rect 161480 4150 161532 4156
rect 160192 3664 160244 3670
rect 160192 3606 160244 3612
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 160204 1850 160232 3606
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 160112 1822 160232 1850
rect 160112 480 160140 1822
rect 161308 480 161336 3470
rect 161400 3398 161428 3470
rect 161388 3392 161440 3398
rect 161388 3334 161440 3340
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 10406
rect 162872 6914 162900 28222
rect 163148 27606 163176 29838
rect 163136 27600 163188 27606
rect 163136 27542 163188 27548
rect 163976 26234 164004 29838
rect 164240 26920 164292 26926
rect 164240 26862 164292 26868
rect 162964 26206 164004 26234
rect 162964 7682 162992 26206
rect 162952 7676 163004 7682
rect 162952 7618 163004 7624
rect 164252 6914 164280 26862
rect 164344 9042 164372 29838
rect 165816 26234 165844 29838
rect 166828 27062 166856 29838
rect 167656 29838 167707 29866
rect 168392 29838 168642 29866
rect 168760 29838 169543 29866
rect 169772 29838 170461 29866
rect 171334 29866 171362 30049
rect 172269 29866 172297 30049
rect 173153 29866 173181 30049
rect 174071 29866 174099 30049
rect 174972 29866 175000 30049
rect 175890 29866 175918 30049
rect 176774 29866 176802 30049
rect 177692 29866 177720 30049
rect 178593 29866 178621 30049
rect 179511 29866 179539 30049
rect 180412 29866 180440 30049
rect 181330 29866 181358 30049
rect 171334 29838 171364 29866
rect 166816 27056 166868 27062
rect 166816 26998 166868 27004
rect 167656 26926 167684 29838
rect 167644 26920 167696 26926
rect 167644 26862 167696 26868
rect 165632 26206 165844 26234
rect 164332 9036 164384 9042
rect 164332 8978 164384 8984
rect 162872 6886 163728 6914
rect 164252 6886 164464 6914
rect 163700 480 163728 6886
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 6886
rect 165632 6186 165660 26206
rect 168392 15978 168420 29838
rect 168760 26234 168788 29838
rect 168484 26206 168788 26234
rect 168484 17338 168512 26206
rect 169772 18698 169800 29838
rect 171336 27606 171364 29838
rect 172256 29838 172297 29866
rect 172532 29838 173181 29866
rect 173912 29838 174099 29866
rect 174924 29838 175000 29866
rect 175844 29838 175918 29866
rect 176764 29838 176802 29866
rect 177684 29838 177720 29866
rect 178052 29838 178621 29866
rect 179432 29838 179539 29866
rect 180352 29838 180440 29866
rect 181272 29838 181358 29866
rect 182231 29866 182259 30049
rect 183149 29866 183177 30049
rect 184050 29866 184078 30049
rect 184968 29866 184996 30049
rect 182231 29838 182312 29866
rect 170404 27600 170456 27606
rect 170404 27542 170456 27548
rect 171324 27600 171376 27606
rect 171324 27542 171376 27548
rect 169760 18692 169812 18698
rect 169760 18634 169812 18640
rect 168472 17332 168524 17338
rect 168472 17274 168524 17280
rect 168380 15972 168432 15978
rect 168380 15914 168432 15920
rect 170312 13184 170364 13190
rect 170312 13126 170364 13132
rect 168380 10668 168432 10674
rect 168380 10610 168432 10616
rect 166080 10600 166132 10606
rect 166080 10542 166132 10548
rect 165620 6180 165672 6186
rect 165620 6122 165672 6128
rect 166092 480 166120 10542
rect 168392 3398 168420 10610
rect 168472 4208 168524 4214
rect 168472 4150 168524 4156
rect 168380 3392 168432 3398
rect 168380 3334 168432 3340
rect 168484 3210 168512 4150
rect 169576 3392 169628 3398
rect 169576 3334 169628 3340
rect 168392 3182 168512 3210
rect 167184 2168 167236 2174
rect 167184 2110 167236 2116
rect 167196 480 167224 2110
rect 168392 480 168420 3182
rect 169588 480 169616 3334
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 13126
rect 170416 4894 170444 27542
rect 172256 26994 172284 29838
rect 172244 26988 172296 26994
rect 172244 26930 172296 26936
rect 172532 20058 172560 29838
rect 173164 27600 173216 27606
rect 173164 27542 173216 27548
rect 172520 20052 172572 20058
rect 172520 19994 172572 20000
rect 172704 10736 172756 10742
rect 172704 10678 172756 10684
rect 170404 4888 170456 4894
rect 170404 4830 170456 4836
rect 171968 4888 172020 4894
rect 171968 4830 172020 4836
rect 171980 480 172008 4830
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 10678
rect 173176 8974 173204 27542
rect 173912 21418 173940 29838
rect 174924 26234 174952 29838
rect 175844 26234 175872 29838
rect 176660 28348 176712 28354
rect 176660 28290 176712 28296
rect 175924 26920 175976 26926
rect 175924 26862 175976 26868
rect 174004 26206 174952 26234
rect 175292 26206 175872 26234
rect 174004 22778 174032 26206
rect 173992 22772 174044 22778
rect 173992 22714 174044 22720
rect 173900 21412 173952 21418
rect 173900 21354 173952 21360
rect 173900 13252 173952 13258
rect 173900 13194 173952 13200
rect 173164 8968 173216 8974
rect 173164 8910 173216 8916
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 13194
rect 175292 5098 175320 26206
rect 175936 7682 175964 26862
rect 175464 7676 175516 7682
rect 175464 7618 175516 7624
rect 175924 7676 175976 7682
rect 175924 7618 175976 7624
rect 175280 5092 175332 5098
rect 175280 5034 175332 5040
rect 175476 480 175504 7618
rect 176672 3874 176700 28290
rect 176764 26926 176792 29838
rect 176752 26920 176804 26926
rect 176752 26862 176804 26868
rect 177684 26234 177712 29838
rect 176764 26206 177712 26234
rect 176764 24138 176792 26206
rect 176752 24132 176804 24138
rect 176752 24074 176804 24080
rect 176752 7812 176804 7818
rect 176752 7754 176804 7760
rect 176660 3868 176712 3874
rect 176660 3810 176712 3816
rect 176764 3482 176792 7754
rect 178052 5370 178080 29838
rect 179052 9036 179104 9042
rect 179052 8978 179104 8984
rect 178040 5364 178092 5370
rect 178040 5306 178092 5312
rect 177856 3868 177908 3874
rect 177856 3810 177908 3816
rect 176672 3454 176792 3482
rect 176672 480 176700 3454
rect 177868 480 177896 3810
rect 179064 480 179092 8978
rect 179432 5030 179460 29838
rect 180352 26234 180380 29838
rect 181272 26234 181300 29838
rect 182180 28144 182232 28150
rect 182180 28086 182232 28092
rect 179524 26206 180380 26234
rect 180812 26206 181300 26234
rect 179420 5024 179472 5030
rect 179420 4966 179472 4972
rect 179524 4962 179552 26206
rect 180812 17270 180840 26206
rect 180800 17264 180852 17270
rect 180800 17206 180852 17212
rect 180248 10804 180300 10810
rect 180248 10746 180300 10752
rect 179512 4956 179564 4962
rect 179512 4898 179564 4904
rect 180260 480 180288 10746
rect 182192 4826 182220 28086
rect 182284 4894 182312 29838
rect 183112 29838 183177 29866
rect 184032 29838 184078 29866
rect 184952 29838 184996 29866
rect 185852 29866 185880 30049
rect 186770 29866 186798 30049
rect 185852 29838 185900 29866
rect 183112 28150 183140 29838
rect 183100 28144 183152 28150
rect 183100 28086 183152 28092
rect 184032 26234 184060 29838
rect 184952 27130 184980 29838
rect 185032 28416 185084 28422
rect 185032 28358 185084 28364
rect 184940 27124 184992 27130
rect 184940 27066 184992 27072
rect 184204 27056 184256 27062
rect 184204 26998 184256 27004
rect 183572 26206 184060 26234
rect 183572 25566 183600 26206
rect 183560 25560 183612 25566
rect 183560 25502 183612 25508
rect 183744 16448 183796 16454
rect 183744 16390 183796 16396
rect 182548 6180 182600 6186
rect 182548 6122 182600 6128
rect 182272 4888 182324 4894
rect 182272 4830 182324 4836
rect 182180 4820 182232 4826
rect 182180 4762 182232 4768
rect 181444 2236 181496 2242
rect 181444 2178 181496 2184
rect 181456 480 181484 2178
rect 182560 480 182588 6122
rect 183756 480 183784 16390
rect 184216 5574 184244 26998
rect 185044 26234 185072 28358
rect 185872 27606 185900 29838
rect 186700 29838 186798 29866
rect 187671 29866 187699 30049
rect 188606 29866 188634 30049
rect 189490 29866 189518 30049
rect 187671 29838 187740 29866
rect 185860 27600 185912 27606
rect 185860 27542 185912 27548
rect 186700 26234 186728 29838
rect 186964 27600 187016 27606
rect 186964 27542 187016 27548
rect 184952 26206 185072 26234
rect 186332 26206 186728 26234
rect 184204 5568 184256 5574
rect 184204 5510 184256 5516
rect 184952 480 184980 26206
rect 186332 19990 186360 26206
rect 186320 19984 186372 19990
rect 186320 19926 186372 19932
rect 186976 18630 187004 27542
rect 186964 18624 187016 18630
rect 186964 18566 187016 18572
rect 187332 7880 187384 7886
rect 187332 7822 187384 7828
rect 186136 5568 186188 5574
rect 186136 5510 186188 5516
rect 186148 480 186176 5510
rect 187344 480 187372 7822
rect 187712 6662 187740 29838
rect 188540 29838 188634 29866
rect 189080 29844 189132 29850
rect 188540 26234 188568 29838
rect 189080 29786 189132 29792
rect 189460 29838 189518 29866
rect 190425 29850 190453 30049
rect 190413 29844 190465 29850
rect 187804 26206 188568 26234
rect 187700 6656 187752 6662
rect 187700 6598 187752 6604
rect 187804 6594 187832 26206
rect 189092 24682 189120 29786
rect 189460 27062 189488 29838
rect 191326 29832 191354 30049
rect 192244 29832 192272 30049
rect 193145 29832 193173 30049
rect 194063 29832 194091 30049
rect 194964 29832 194992 30049
rect 195882 29832 195910 30049
rect 190413 29786 190465 29792
rect 191024 29804 191354 29832
rect 191852 29804 192272 29832
rect 193140 29804 193173 29832
rect 193232 29804 194091 29832
rect 194704 29804 194992 29832
rect 195808 29804 195910 29832
rect 196783 29832 196811 30049
rect 197452 29844 197504 29850
rect 196783 29804 196848 29832
rect 189448 27056 189500 27062
rect 189448 26998 189500 27004
rect 191024 26234 191052 29804
rect 191104 26988 191156 26994
rect 191104 26930 191156 26936
rect 190472 26206 191052 26234
rect 189080 24676 189132 24682
rect 189080 24618 189132 24624
rect 188528 11756 188580 11762
rect 188528 11698 188580 11704
rect 187792 6588 187844 6594
rect 187792 6530 187844 6536
rect 188540 480 188568 11698
rect 189724 7676 189776 7682
rect 189724 7618 189776 7624
rect 189736 480 189764 7618
rect 190472 6526 190500 26206
rect 190828 9376 190880 9382
rect 190828 9318 190880 9324
rect 190460 6520 190512 6526
rect 190460 6462 190512 6468
rect 190840 480 190868 9318
rect 191116 7682 191144 26930
rect 191104 7676 191156 7682
rect 191104 7618 191156 7624
rect 191852 6458 191880 29804
rect 193140 26994 193168 29804
rect 191932 26988 191984 26994
rect 191932 26930 191984 26936
rect 193128 26988 193180 26994
rect 193128 26930 193180 26936
rect 191840 6452 191892 6458
rect 191840 6394 191892 6400
rect 191944 6390 191972 26930
rect 191932 6384 191984 6390
rect 191932 6326 191984 6332
rect 193232 6322 193260 29804
rect 194600 28484 194652 28490
rect 194600 28426 194652 28432
rect 193312 22024 193364 22030
rect 193312 21966 193364 21972
rect 193220 6316 193272 6322
rect 193220 6258 193272 6264
rect 193220 3868 193272 3874
rect 193220 3810 193272 3816
rect 192024 2304 192076 2310
rect 192024 2246 192076 2252
rect 192036 480 192064 2246
rect 193232 480 193260 3810
rect 193324 3482 193352 21966
rect 193404 15972 193456 15978
rect 193404 15914 193456 15920
rect 193416 3874 193444 15914
rect 193404 3868 193456 3874
rect 193404 3810 193456 3816
rect 193324 3454 194456 3482
rect 194428 480 194456 3454
rect 194612 490 194640 28426
rect 194704 6254 194732 29804
rect 195808 26234 195836 29804
rect 196820 27198 196848 29804
rect 197684 29832 197712 30049
rect 198585 29850 198613 30049
rect 197452 29786 197504 29792
rect 197648 29804 197712 29832
rect 198573 29844 198625 29850
rect 196808 27192 196860 27198
rect 196808 27134 196860 27140
rect 194796 26206 195836 26234
rect 194692 6248 194744 6254
rect 194692 6190 194744 6196
rect 194796 6186 194824 26206
rect 197360 25968 197412 25974
rect 197360 25910 197412 25916
rect 195980 17332 196032 17338
rect 195980 17274 196032 17280
rect 195992 16574 196020 17274
rect 197372 16574 197400 25910
rect 197464 21962 197492 29786
rect 197648 26234 197676 29804
rect 199503 29832 199531 30049
rect 198573 29786 198625 29792
rect 198752 29804 199531 29832
rect 200120 29844 200172 29850
rect 197556 26206 197676 26234
rect 197556 23322 197584 26206
rect 198752 24614 198780 29804
rect 200421 29832 200449 30049
rect 201322 29850 201350 30049
rect 200120 29786 200172 29792
rect 200224 29804 200449 29832
rect 201310 29844 201362 29850
rect 199384 27056 199436 27062
rect 199384 26998 199436 27004
rect 198740 24608 198792 24614
rect 198740 24550 198792 24556
rect 197544 23316 197596 23322
rect 197544 23258 197596 23264
rect 197452 21956 197504 21962
rect 197452 21898 197504 21904
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194784 6180 194836 6186
rect 194784 6122 194836 6128
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 194612 462 195192 490
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 199396 8022 199424 26998
rect 199384 8016 199436 8022
rect 199384 7958 199436 7964
rect 200132 7750 200160 29786
rect 200224 26042 200252 29804
rect 202240 29832 202268 30049
rect 201310 29786 201362 29792
rect 202156 29804 202268 29832
rect 203158 29832 203186 30049
rect 204059 29832 204087 30049
rect 204977 29832 205005 30049
rect 203158 29804 203196 29832
rect 204059 29804 204116 29832
rect 201500 28552 201552 28558
rect 201500 28494 201552 28500
rect 200212 26036 200264 26042
rect 200212 25978 200264 25984
rect 200212 18692 200264 18698
rect 200212 18634 200264 18640
rect 200224 16574 200252 18634
rect 200224 16546 200344 16574
rect 200120 7744 200172 7750
rect 200120 7686 200172 7692
rect 199108 2372 199160 2378
rect 199108 2314 199160 2320
rect 199120 480 199148 2314
rect 200316 480 200344 16546
rect 201512 3398 201540 28494
rect 202156 26234 202184 29804
rect 203168 27334 203196 29804
rect 204088 27606 204116 29804
rect 204272 29804 205005 29832
rect 205640 29844 205692 29850
rect 204076 27600 204128 27606
rect 204076 27542 204128 27548
rect 203156 27328 203208 27334
rect 203156 27270 203208 27276
rect 201604 26206 202184 26234
rect 201604 17746 201632 26206
rect 204272 19038 204300 29804
rect 205878 29832 205906 30049
rect 206762 29850 206790 30049
rect 205640 29786 205692 29792
rect 205836 29804 205906 29832
rect 206750 29844 206802 29850
rect 205548 27600 205600 27606
rect 205548 27542 205600 27548
rect 205560 20466 205588 27542
rect 205652 23254 205680 29786
rect 205836 26234 205864 29804
rect 207697 29832 207725 30049
rect 208598 29832 208626 30049
rect 209499 29832 209527 30049
rect 210451 29832 210479 30049
rect 206750 29786 206802 29792
rect 207676 29804 207725 29832
rect 208412 29804 208626 29832
rect 208688 29804 209527 29832
rect 209792 29804 210479 29832
rect 211160 29844 211212 29850
rect 207676 27402 207704 29804
rect 207664 27396 207716 27402
rect 207664 27338 207716 27344
rect 205744 26206 205864 26234
rect 205744 24478 205772 26206
rect 205732 24472 205784 24478
rect 205732 24414 205784 24420
rect 205640 23248 205692 23254
rect 205640 23190 205692 23196
rect 208412 21690 208440 29804
rect 208688 26234 208716 29804
rect 208504 26206 208716 26234
rect 208504 25906 208532 26206
rect 208492 25900 208544 25906
rect 208492 25842 208544 25848
rect 208400 21684 208452 21690
rect 208400 21626 208452 21632
rect 205548 20460 205600 20466
rect 205548 20402 205600 20408
rect 204260 19032 204312 19038
rect 204260 18974 204312 18980
rect 201592 17740 201644 17746
rect 201592 17682 201644 17688
rect 208584 16516 208636 16522
rect 208584 16458 208636 16464
rect 206192 14544 206244 14550
rect 206192 14486 206244 14492
rect 203892 8968 203944 8974
rect 203892 8910 203944 8916
rect 201592 5296 201644 5302
rect 201592 5238 201644 5244
rect 201500 3392 201552 3398
rect 201500 3334 201552 3340
rect 201604 2666 201632 5238
rect 202696 3392 202748 3398
rect 202696 3334 202748 3340
rect 201512 2638 201632 2666
rect 201512 480 201540 2638
rect 202708 480 202736 3334
rect 203904 480 203932 8910
rect 205088 7948 205140 7954
rect 205088 7890 205140 7896
rect 205100 480 205128 7890
rect 206204 480 206232 14486
rect 207388 7676 207440 7682
rect 207388 7618 207440 7624
rect 207400 480 207428 7618
rect 208596 480 208624 16458
rect 209792 7682 209820 29804
rect 211318 29832 211346 30049
rect 212253 29850 212281 30049
rect 211160 29786 211212 29792
rect 211264 29804 211346 29832
rect 212241 29844 212293 29850
rect 211172 20330 211200 29786
rect 211160 20324 211212 20330
rect 211160 20266 211212 20272
rect 209872 20052 209924 20058
rect 209872 19994 209924 20000
rect 209780 7676 209832 7682
rect 209780 7618 209832 7624
rect 209884 3874 209912 19994
rect 211160 17808 211212 17814
rect 211160 17750 211212 17756
rect 211172 16574 211200 17750
rect 211264 17678 211292 29804
rect 213137 29832 213165 30049
rect 214072 29832 214100 30049
rect 214973 29832 215001 30049
rect 215891 29832 215919 30049
rect 216792 29832 216820 30049
rect 217727 29832 217755 30049
rect 218577 29832 218605 30049
rect 212241 29786 212293 29792
rect 212552 29804 213165 29832
rect 214024 29804 214100 29832
rect 214944 29804 215001 29832
rect 215312 29804 215919 29832
rect 216692 29804 216820 29832
rect 216968 29804 217755 29832
rect 218164 29804 218605 29832
rect 212552 18970 212580 29804
rect 214024 26234 214052 29804
rect 214944 27470 214972 29804
rect 214932 27464 214984 27470
rect 214932 27406 214984 27412
rect 213932 26206 214052 26234
rect 213932 24410 213960 26206
rect 213920 24404 213972 24410
rect 213920 24346 213972 24352
rect 215312 23118 215340 29804
rect 215300 23112 215352 23118
rect 215300 23054 215352 23060
rect 216692 21758 216720 29804
rect 216968 26234 216996 29804
rect 216784 26206 216996 26234
rect 216784 25838 216812 26206
rect 216772 25832 216824 25838
rect 216772 25774 216824 25780
rect 218060 22772 218112 22778
rect 218060 22714 218112 22720
rect 216680 21752 216732 21758
rect 216680 21694 216732 21700
rect 213920 21412 213972 21418
rect 213920 21354 213972 21360
rect 212540 18964 212592 18970
rect 212540 18906 212592 18912
rect 211252 17672 211304 17678
rect 211252 17614 211304 17620
rect 213932 16574 213960 21354
rect 211172 16546 211752 16574
rect 213932 16546 214512 16574
rect 209964 14612 210016 14618
rect 209964 14554 210016 14560
rect 209872 3868 209924 3874
rect 209872 3810 209924 3816
rect 209976 3482 210004 14554
rect 210976 3868 211028 3874
rect 210976 3810 211028 3816
rect 209792 3454 210004 3482
rect 209792 480 209820 3454
rect 210988 480 211016 3810
rect 195164 354 195192 462
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213368 14680 213420 14686
rect 213368 14622 213420 14628
rect 213380 480 213408 14622
rect 214484 480 214512 16546
rect 216864 14748 216916 14754
rect 216864 14690 216916 14696
rect 215300 11892 215352 11898
rect 215300 11834 215352 11840
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 11834
rect 216876 480 216904 14690
rect 218072 480 218100 22714
rect 218164 17610 218192 29804
rect 219529 29730 219557 30049
rect 220413 29866 220441 30049
rect 221331 29866 221359 30049
rect 219728 29838 220441 29866
rect 220832 29838 221359 29866
rect 222249 29866 222277 30049
rect 223150 29866 223178 30049
rect 224068 29866 224096 30049
rect 222249 29838 222332 29866
rect 219529 29702 219572 29730
rect 219544 27266 219572 29702
rect 219532 27260 219584 27266
rect 219532 27202 219584 27208
rect 219728 26234 219756 29838
rect 219452 26206 219756 26234
rect 219452 20262 219480 26206
rect 219440 20256 219492 20262
rect 219440 20198 219492 20204
rect 220832 18902 220860 29838
rect 222200 28144 222252 28150
rect 222200 28086 222252 28092
rect 220820 18896 220872 18902
rect 220820 18838 220872 18844
rect 218152 17604 218204 17610
rect 218152 17546 218204 17552
rect 219992 14816 220044 14822
rect 219992 14758 220044 14764
rect 219256 11960 219308 11966
rect 219256 11902 219308 11908
rect 219268 480 219296 11902
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 14758
rect 222212 9246 222240 28086
rect 222304 9314 222332 29838
rect 223132 29838 223178 29866
rect 224052 29838 224096 29866
rect 224969 29866 224997 30049
rect 225887 29866 225915 30049
rect 226805 29866 226833 30049
rect 224969 29838 225000 29866
rect 225887 29838 225920 29866
rect 223132 28150 223160 29838
rect 223120 28144 223172 28150
rect 223120 28086 223172 28092
rect 224052 26234 224080 29838
rect 224224 26920 224276 26926
rect 224224 26862 224276 26868
rect 223592 26206 224080 26234
rect 222752 12028 222804 12034
rect 222752 11970 222804 11976
rect 222292 9308 222344 9314
rect 222292 9250 222344 9256
rect 222200 9240 222252 9246
rect 222200 9182 222252 9188
rect 221556 5092 221608 5098
rect 221556 5034 221608 5040
rect 221568 480 221596 5034
rect 222764 480 222792 11970
rect 223592 9178 223620 26206
rect 223580 9172 223632 9178
rect 223580 9114 223632 9120
rect 224236 8294 224264 26862
rect 224972 24342 225000 29838
rect 225892 27538 225920 29838
rect 226352 29838 226833 29866
rect 227706 29866 227734 30049
rect 228624 29866 228652 30049
rect 229542 29866 229570 30049
rect 230409 29866 230437 30049
rect 231344 29866 231372 30049
rect 232245 29866 232273 30049
rect 227706 29838 227760 29866
rect 225880 27532 225932 27538
rect 225880 27474 225932 27480
rect 224960 24336 225012 24342
rect 224960 24278 225012 24284
rect 226352 9110 226380 29838
rect 227732 26234 227760 29838
rect 228560 29838 228652 29866
rect 229480 29838 229570 29866
rect 230400 29838 230437 29866
rect 231320 29838 231372 29866
rect 231860 29844 231912 29850
rect 228560 26234 228588 29838
rect 229480 26234 229508 29838
rect 230400 26926 230428 29838
rect 230388 26920 230440 26926
rect 230388 26862 230440 26868
rect 231320 26234 231348 29838
rect 231860 29786 231912 29792
rect 231964 29838 232273 29866
rect 233146 29850 233174 30049
rect 234081 29866 234109 30049
rect 234965 29866 234993 30049
rect 235900 29866 235928 30049
rect 236801 29866 236829 30049
rect 237719 29866 237747 30049
rect 233134 29844 233186 29850
rect 227732 26206 227852 26234
rect 227720 24132 227772 24138
rect 227720 24074 227772 24080
rect 226432 17536 226484 17542
rect 226432 17478 226484 17484
rect 226340 9104 226392 9110
rect 226340 9046 226392 9052
rect 224224 8288 224276 8294
rect 224224 8230 224276 8236
rect 225144 8288 225196 8294
rect 225144 8230 225196 8236
rect 223948 5228 224000 5234
rect 223948 5170 224000 5176
rect 223960 480 223988 5170
rect 225156 480 225184 8230
rect 226444 3874 226472 17478
rect 226524 12096 226576 12102
rect 226524 12038 226576 12044
rect 226432 3868 226484 3874
rect 226432 3810 226484 3816
rect 226536 3482 226564 12038
rect 227732 6914 227760 24074
rect 227824 9042 227852 26206
rect 227916 26206 228588 26234
rect 229112 26206 229508 26234
rect 230492 26206 231348 26234
rect 227916 22982 227944 26206
rect 227904 22976 227956 22982
rect 227904 22918 227956 22924
rect 229112 21622 229140 26206
rect 229100 21616 229152 21622
rect 229100 21558 229152 21564
rect 229376 10872 229428 10878
rect 229376 10814 229428 10820
rect 227812 9036 227864 9042
rect 227812 8978 227864 8984
rect 227732 6886 228312 6914
rect 227536 3868 227588 3874
rect 227536 3810 227588 3816
rect 226352 3454 226564 3482
rect 226352 480 226380 3454
rect 227548 480 227576 3810
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 6886
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 10814
rect 230492 8974 230520 26206
rect 231032 14952 231084 14958
rect 231032 14894 231084 14900
rect 230480 8968 230532 8974
rect 230480 8910 230532 8916
rect 231044 480 231072 14894
rect 231872 5166 231900 29786
rect 231964 25770 231992 29838
rect 233134 29786 233186 29792
rect 233252 29838 234109 29866
rect 234632 29838 234993 29866
rect 235828 29838 235928 29866
rect 236012 29838 236829 29866
rect 237380 29844 237432 29850
rect 231952 25764 232004 25770
rect 231952 25706 232004 25712
rect 233252 17474 233280 29838
rect 233240 17468 233292 17474
rect 233240 17410 233292 17416
rect 234632 13326 234660 29838
rect 235828 26234 235856 29838
rect 234724 26206 235856 26234
rect 234724 20194 234752 26206
rect 236012 24274 236040 29838
rect 237380 29786 237432 29792
rect 237484 29838 237747 29866
rect 238620 29850 238648 30049
rect 238608 29844 238660 29850
rect 236000 24268 236052 24274
rect 236000 24210 236052 24216
rect 234712 20188 234764 20194
rect 234712 20130 234764 20136
rect 234620 13320 234672 13326
rect 234620 13262 234672 13268
rect 236552 12232 236604 12238
rect 236552 12174 236604 12180
rect 233424 12164 233476 12170
rect 233424 12106 233476 12112
rect 232228 5364 232280 5370
rect 232228 5306 232280 5312
rect 231860 5160 231912 5166
rect 231860 5102 231912 5108
rect 232240 480 232268 5306
rect 233436 480 233464 12106
rect 235816 5024 235868 5030
rect 235816 4966 235868 4972
rect 234620 3868 234672 3874
rect 234620 3810 234672 3816
rect 234632 480 234660 3810
rect 235828 480 235856 4966
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 12174
rect 237392 2106 237420 29786
rect 237484 18834 237512 29838
rect 239538 29832 239566 30049
rect 238608 29786 238660 29792
rect 239508 29804 239566 29832
rect 240140 29844 240192 29850
rect 239508 26234 239536 29804
rect 240439 29832 240467 30049
rect 241374 29850 241402 30049
rect 242224 29866 242252 30049
rect 240140 29786 240192 29792
rect 240428 29804 240467 29832
rect 241362 29844 241414 29850
rect 238772 26206 239536 26234
rect 237472 18828 237524 18834
rect 237472 18770 237524 18776
rect 237656 15972 237708 15978
rect 237656 15914 237708 15920
rect 237380 2100 237432 2106
rect 237380 2042 237432 2048
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 15914
rect 238772 10402 238800 26206
rect 238760 10396 238812 10402
rect 238760 10338 238812 10344
rect 240152 10334 240180 29786
rect 240428 27062 240456 29804
rect 242224 29838 242296 29866
rect 241362 29786 241414 29792
rect 242164 27192 242216 27198
rect 242164 27134 242216 27140
rect 240416 27056 240468 27062
rect 240416 26998 240468 27004
rect 241704 16040 241756 16046
rect 241704 15982 241756 15988
rect 240140 10328 240192 10334
rect 240140 10270 240192 10276
rect 240508 5364 240560 5370
rect 240508 5306 240560 5312
rect 239312 4956 239364 4962
rect 239312 4898 239364 4904
rect 239324 480 239352 4898
rect 240520 480 240548 5306
rect 241716 480 241744 15982
rect 242176 8090 242204 27134
rect 242268 26994 242296 29838
rect 242900 29844 242952 29850
rect 243159 29832 243187 30049
rect 244060 29850 244088 30049
rect 244048 29844 244100 29850
rect 243159 29804 243216 29832
rect 242900 29786 242952 29792
rect 242256 26988 242308 26994
rect 242256 26930 242308 26936
rect 242912 18766 242940 29786
rect 243188 27606 243216 29804
rect 244978 29832 245006 30049
rect 245896 29832 245924 30049
rect 246797 29832 246825 30049
rect 247715 29832 247743 30049
rect 248633 29866 248661 30049
rect 244048 29786 244100 29792
rect 244936 29804 245006 29832
rect 245672 29804 245924 29832
rect 246040 29804 246825 29832
rect 247052 29804 247743 29832
rect 248432 29838 248661 29866
rect 249534 29866 249562 30049
rect 250452 29866 250480 30049
rect 251353 29866 251381 30049
rect 252271 29866 252299 30049
rect 253189 29866 253217 30049
rect 254056 29866 254084 30049
rect 254974 29866 255002 30049
rect 255892 29866 255920 30049
rect 256793 29866 256821 30049
rect 257728 29866 257756 30049
rect 249534 29838 249564 29866
rect 244936 29594 244964 29804
rect 244844 29566 244964 29594
rect 243176 27600 243228 27606
rect 243176 27542 243228 27548
rect 244844 26234 244872 29566
rect 244924 27600 244976 27606
rect 244924 27542 244976 27548
rect 244292 26206 244872 26234
rect 244292 21554 244320 26206
rect 244280 21548 244332 21554
rect 244280 21490 244332 21496
rect 242900 18760 242952 18766
rect 242900 18702 242952 18708
rect 244936 17406 244964 27542
rect 245672 20126 245700 29804
rect 246040 26234 246068 29804
rect 246304 27124 246356 27130
rect 246304 27066 246356 27072
rect 245764 26206 246068 26234
rect 245764 22914 245792 26206
rect 245752 22908 245804 22914
rect 245752 22850 245804 22856
rect 245660 20120 245712 20126
rect 245660 20062 245712 20068
rect 244924 17400 244976 17406
rect 244924 17342 244976 17348
rect 242900 17264 242952 17270
rect 242900 17206 242952 17212
rect 242164 8084 242216 8090
rect 242164 8026 242216 8032
rect 242912 480 242940 17206
rect 245200 16176 245252 16182
rect 245200 16118 245252 16124
rect 244096 8220 244148 8226
rect 244096 8162 244148 8168
rect 244108 480 244136 8162
rect 245212 480 245240 16118
rect 246316 5438 246344 27066
rect 247052 25702 247080 29804
rect 247040 25696 247092 25702
rect 247040 25638 247092 25644
rect 248432 24206 248460 29838
rect 249064 27532 249116 27538
rect 249064 27474 249116 27480
rect 248420 24200 248472 24206
rect 248420 24142 248472 24148
rect 248420 16244 248472 16250
rect 248420 16186 248472 16192
rect 247592 12300 247644 12306
rect 247592 12242 247644 12248
rect 246304 5432 246356 5438
rect 246304 5374 246356 5380
rect 246396 4888 246448 4894
rect 246396 4830 246448 4836
rect 246408 480 246436 4830
rect 247604 480 247632 12242
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 16186
rect 249076 13394 249104 27474
rect 249536 27130 249564 29838
rect 250364 29838 250480 29866
rect 251284 29838 251381 29866
rect 251652 29838 252299 29866
rect 252664 29838 253217 29866
rect 254044 29838 254084 29866
rect 254964 29838 255002 29866
rect 255884 29838 255920 29866
rect 256712 29838 256821 29866
rect 257724 29838 257756 29866
rect 249524 27124 249576 27130
rect 249524 27066 249576 27072
rect 250364 26234 250392 29838
rect 249812 26206 250392 26234
rect 249064 13388 249116 13394
rect 249064 13330 249116 13336
rect 249812 5098 249840 26206
rect 251180 21820 251232 21826
rect 251180 21762 251232 21768
rect 249800 5092 249852 5098
rect 249800 5034 249852 5040
rect 249984 4820 250036 4826
rect 249984 4762 250036 4768
rect 249996 480 250024 4762
rect 251192 3942 251220 21762
rect 251284 17338 251312 29838
rect 251652 26234 251680 29838
rect 251376 26206 251680 26234
rect 251376 18698 251404 26206
rect 252560 25560 252612 25566
rect 252560 25502 252612 25508
rect 251364 18692 251416 18698
rect 251364 18634 251416 18640
rect 251272 17332 251324 17338
rect 251272 17274 251324 17280
rect 252572 16574 252600 25502
rect 252664 21486 252692 29838
rect 254044 27606 254072 29838
rect 254032 27600 254084 27606
rect 254032 27542 254084 27548
rect 254964 26234 254992 29838
rect 255884 26234 255912 29838
rect 256608 27600 256660 27606
rect 256608 27542 256660 27548
rect 253952 26206 254992 26234
rect 255332 26206 255912 26234
rect 253952 22846 253980 26206
rect 253940 22840 253992 22846
rect 253940 22782 253992 22788
rect 252652 21480 252704 21486
rect 252652 21422 252704 21428
rect 252572 16546 253520 16574
rect 251272 10940 251324 10946
rect 251272 10882 251324 10888
rect 251180 3936 251232 3942
rect 251180 3878 251232 3884
rect 251284 3482 251312 10882
rect 252376 3936 252428 3942
rect 252376 3878 252428 3884
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3878
rect 253492 480 253520 16546
rect 254676 9512 254728 9518
rect 254676 9454 254728 9460
rect 254688 480 254716 9454
rect 255332 5030 255360 26206
rect 256620 20058 256648 27542
rect 256608 20052 256660 20058
rect 256608 19994 256660 20000
rect 255872 16312 255924 16318
rect 255872 16254 255924 16260
rect 255320 5024 255372 5030
rect 255320 4966 255372 4972
rect 255884 480 255912 16254
rect 256712 4962 256740 29838
rect 257724 26234 257752 29838
rect 258612 29832 258640 30049
rect 258552 29804 258640 29832
rect 259460 29844 259512 29850
rect 258552 26234 258580 29804
rect 259547 29832 259575 30049
rect 260448 29850 260476 30049
rect 260436 29844 260488 29850
rect 259547 29804 259592 29832
rect 259460 29786 259512 29792
rect 256804 26206 257752 26234
rect 258092 26206 258580 26234
rect 256700 4956 256752 4962
rect 256700 4898 256752 4904
rect 256804 4894 256832 26206
rect 257068 5432 257120 5438
rect 257068 5374 257120 5380
rect 256792 4888 256844 4894
rect 256792 4830 256844 4836
rect 257080 480 257108 5374
rect 258092 4826 258120 26206
rect 259472 24138 259500 29786
rect 259564 25634 259592 29804
rect 261366 29832 261394 30049
rect 262267 29832 262295 30049
rect 263202 29832 263230 30049
rect 264086 29832 264114 30049
rect 265021 29832 265049 30049
rect 265871 29832 265899 30049
rect 266806 29832 266834 30049
rect 261366 29804 261432 29832
rect 260436 29786 260488 29792
rect 261404 27198 261432 29804
rect 262232 29804 262295 29832
rect 263152 29804 263230 29832
rect 264072 29804 264114 29832
rect 264992 29804 265049 29832
rect 265176 29804 265899 29832
rect 266740 29804 266834 29832
rect 267707 29832 267735 30049
rect 268625 29832 268653 30049
rect 269543 29832 269571 30049
rect 270444 29832 270472 30049
rect 271362 29832 271390 30049
rect 272280 29832 272308 30049
rect 273181 29832 273209 30049
rect 274099 29832 274127 30049
rect 267707 29804 267780 29832
rect 261392 27192 261444 27198
rect 261392 27134 261444 27140
rect 259552 25628 259604 25634
rect 259552 25570 259604 25576
rect 259460 24132 259512 24138
rect 259460 24074 259512 24080
rect 259460 18624 259512 18630
rect 259460 18566 259512 18572
rect 259472 11694 259500 18566
rect 262232 17270 262260 29804
rect 263152 26234 263180 29804
rect 264072 26234 264100 29804
rect 264992 27606 265020 29804
rect 264980 27600 265032 27606
rect 264980 27542 265032 27548
rect 265176 26234 265204 29804
rect 266740 26234 266768 29804
rect 267648 27600 267700 27606
rect 267648 27542 267700 27548
rect 262324 26206 263180 26234
rect 263612 26206 264100 26234
rect 264992 26206 265204 26234
rect 266372 26206 266768 26234
rect 262324 18630 262352 26206
rect 263612 21418 263640 26206
rect 264992 22778 265020 26206
rect 266372 25566 266400 26206
rect 266360 25560 266412 25566
rect 266360 25502 266412 25508
rect 264980 22772 265032 22778
rect 264980 22714 265032 22720
rect 263600 21412 263652 21418
rect 263600 21354 263652 21360
rect 267660 19990 267688 27542
rect 263600 19984 263652 19990
rect 263600 19926 263652 19932
rect 267648 19984 267700 19990
rect 267648 19926 267700 19932
rect 262312 18624 262364 18630
rect 262312 18566 262364 18572
rect 262220 17264 262272 17270
rect 262220 17206 262272 17212
rect 263612 16574 263640 19926
rect 263612 16546 264192 16574
rect 259552 16380 259604 16386
rect 259552 16322 259604 16328
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 258264 8288 258316 8294
rect 258264 8230 258316 8236
rect 258080 4820 258132 4826
rect 258080 4762 258132 4768
rect 258276 480 258304 8230
rect 259564 6914 259592 16322
rect 261760 12368 261812 12374
rect 261760 12310 261812 12316
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 12310
rect 262956 3936 263008 3942
rect 262956 3878 263008 3884
rect 262968 480 262996 3878
rect 264164 480 264192 16546
rect 267752 16114 267780 29804
rect 267844 29804 268653 29832
rect 269132 29804 269571 29832
rect 270420 29804 270472 29832
rect 271340 29804 271390 29832
rect 271892 29804 272308 29832
rect 273180 29804 273209 29832
rect 273364 29804 274127 29832
rect 274640 29844 274692 29850
rect 267844 23050 267872 29804
rect 267832 23044 267884 23050
rect 267832 22986 267884 22992
rect 267740 16108 267792 16114
rect 267740 16050 267792 16056
rect 268384 13728 268436 13734
rect 268384 13670 268436 13676
rect 264980 11008 265032 11014
rect 264980 10950 265032 10956
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 10950
rect 266544 6724 266596 6730
rect 266544 6666 266596 6672
rect 266556 480 266584 6666
rect 267740 6656 267792 6662
rect 267740 6598 267792 6604
rect 267752 480 267780 6598
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 13670
rect 269132 11830 269160 29804
rect 270420 28150 270448 29804
rect 269212 28144 269264 28150
rect 269212 28086 269264 28092
rect 270408 28144 270460 28150
rect 270408 28086 270460 28092
rect 269224 20398 269252 28086
rect 271340 26234 271368 29804
rect 270512 26206 271368 26234
rect 269212 20392 269264 20398
rect 269212 20334 269264 20340
rect 270512 19106 270540 26206
rect 271892 21894 271920 29804
rect 273180 26858 273208 29804
rect 271972 26852 272024 26858
rect 271972 26794 272024 26800
rect 273168 26852 273220 26858
rect 273168 26794 273220 26800
rect 271984 23186 272012 26794
rect 271972 23180 272024 23186
rect 271972 23122 272024 23128
rect 273260 23180 273312 23186
rect 273260 23122 273312 23128
rect 271880 21888 271932 21894
rect 271880 21830 271932 21836
rect 270500 19100 270552 19106
rect 270500 19042 270552 19048
rect 269120 11824 269172 11830
rect 269120 11766 269172 11772
rect 269764 10532 269816 10538
rect 269764 10474 269816 10480
rect 269776 3874 269804 10474
rect 271236 6588 271288 6594
rect 271236 6530 271288 6536
rect 272432 6588 272484 6594
rect 272432 6530 272484 6536
rect 269764 3868 269816 3874
rect 269764 3810 269816 3816
rect 270040 3392 270092 3398
rect 270040 3334 270092 3340
rect 270052 480 270080 3334
rect 271248 480 271276 6530
rect 272444 480 272472 6530
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 23122
rect 273364 13462 273392 29804
rect 275017 29832 275045 30049
rect 275901 29850 275929 30049
rect 274640 29786 274692 29792
rect 274744 29804 275045 29832
rect 275889 29844 275941 29850
rect 273904 27464 273956 27470
rect 273904 27406 273956 27412
rect 273916 13666 273944 27406
rect 273904 13660 273956 13666
rect 273904 13602 273956 13608
rect 274652 13598 274680 29786
rect 274640 13592 274692 13598
rect 274640 13534 274692 13540
rect 274744 13530 274772 29804
rect 276836 29832 276864 30049
rect 277703 29866 277731 30049
rect 275889 29786 275941 29792
rect 276768 29804 276864 29832
rect 277492 29844 277544 29850
rect 276768 26234 276796 29804
rect 277492 29786 277544 29792
rect 277596 29838 277731 29866
rect 278621 29850 278649 30049
rect 279539 29866 279567 30049
rect 280440 29866 280468 30049
rect 281375 29866 281403 30049
rect 282276 29866 282304 30049
rect 278609 29844 278661 29850
rect 276032 26206 276796 26234
rect 274732 13524 274784 13530
rect 274732 13466 274784 13472
rect 273352 13456 273404 13462
rect 273352 13398 273404 13404
rect 273904 11824 273956 11830
rect 273904 11766 273956 11772
rect 273916 3942 273944 11766
rect 276032 10470 276060 26206
rect 277400 24676 277452 24682
rect 277400 24618 277452 24624
rect 276664 24540 276716 24546
rect 276664 24482 276716 24488
rect 276020 10464 276072 10470
rect 276020 10406 276072 10412
rect 274824 8016 274876 8022
rect 274824 7958 274876 7964
rect 273904 3936 273956 3942
rect 273904 3878 273956 3884
rect 274836 480 274864 7958
rect 276020 6656 276072 6662
rect 276020 6598 276072 6604
rect 276032 480 276060 6598
rect 276676 3398 276704 24482
rect 277412 6914 277440 24618
rect 277504 10674 277532 29786
rect 277492 10668 277544 10674
rect 277492 10610 277544 10616
rect 277596 10606 277624 29838
rect 278609 29786 278661 29792
rect 278792 29838 279567 29866
rect 280172 29838 280468 29866
rect 280632 29838 281403 29866
rect 282104 29838 282304 29866
rect 278792 10742 278820 29838
rect 278780 10736 278832 10742
rect 278780 10678 278832 10684
rect 277584 10600 277636 10606
rect 277584 10542 277636 10548
rect 280172 7818 280200 29838
rect 280632 26234 280660 29838
rect 282104 26234 282132 29838
rect 283194 29730 283222 30049
rect 284095 29866 284123 30049
rect 285013 29866 285041 30049
rect 285914 29866 285942 30049
rect 283392 29838 284123 29866
rect 284312 29838 285041 29866
rect 285680 29844 285732 29850
rect 283194 29702 283236 29730
rect 283208 27606 283236 29702
rect 282184 27600 282236 27606
rect 282184 27542 282236 27548
rect 283196 27600 283248 27606
rect 283196 27542 283248 27548
rect 280264 26206 280660 26234
rect 281552 26206 282132 26234
rect 280264 10810 280292 26206
rect 281552 16454 281580 26206
rect 281540 16448 281592 16454
rect 281540 16390 281592 16396
rect 280252 10804 280304 10810
rect 280252 10746 280304 10752
rect 282092 8152 282144 8158
rect 282092 8094 282144 8100
rect 280160 7812 280212 7818
rect 280160 7754 280212 7760
rect 277412 6886 278360 6914
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 276664 3392 276716 3398
rect 276664 3334 276716 3340
rect 277136 480 277164 3810
rect 278332 480 278360 6886
rect 279516 6860 279568 6866
rect 279516 6802 279568 6808
rect 279528 480 279556 6802
rect 281908 6520 281960 6526
rect 281908 6462 281960 6468
rect 280712 3188 280764 3194
rect 280712 3130 280764 3136
rect 280724 480 280752 3130
rect 281920 480 281948 6462
rect 282104 3874 282132 8094
rect 282196 7886 282224 27542
rect 283392 26234 283420 29838
rect 283116 26206 283420 26234
rect 283116 16574 283144 26206
rect 284312 22030 284340 29838
rect 285680 29786 285732 29792
rect 285876 29838 285942 29866
rect 286849 29850 286877 30049
rect 286837 29844 286889 29850
rect 284300 22024 284352 22030
rect 284300 21966 284352 21972
rect 284300 20392 284352 20398
rect 284300 20334 284352 20340
rect 283024 16546 283144 16574
rect 283024 9382 283052 16546
rect 283104 10464 283156 10470
rect 283104 10406 283156 10412
rect 283012 9376 283064 9382
rect 283012 9318 283064 9324
rect 282184 7880 282236 7886
rect 282184 7822 282236 7828
rect 282092 3868 282144 3874
rect 282092 3810 282144 3816
rect 283116 480 283144 10406
rect 284312 480 284340 20334
rect 284944 13524 284996 13530
rect 284944 13466 284996 13472
rect 284956 3194 284984 13466
rect 285404 6452 285456 6458
rect 285404 6394 285456 6400
rect 284944 3188 284996 3194
rect 284944 3130 284996 3136
rect 285416 480 285444 6394
rect 285692 5302 285720 29786
rect 285876 26234 285904 29838
rect 286837 29786 286889 29792
rect 287716 26234 287744 30049
rect 288668 29832 288696 30049
rect 289518 29832 289546 30049
rect 290453 29832 290481 30049
rect 285784 26206 285904 26234
rect 287072 26206 287744 26234
rect 288452 29804 288696 29832
rect 289464 29804 289546 29832
rect 289832 29804 290481 29832
rect 291200 29844 291252 29850
rect 285784 25974 285812 26206
rect 285772 25968 285824 25974
rect 285772 25910 285824 25916
rect 287072 7954 287100 26206
rect 288452 16522 288480 29804
rect 289464 26234 289492 29804
rect 288544 26206 289492 26234
rect 288544 17814 288572 26206
rect 288532 17808 288584 17814
rect 288532 17750 288584 17756
rect 288440 16516 288492 16522
rect 288440 16458 288492 16464
rect 289832 11898 289860 29804
rect 291354 29832 291382 30049
rect 292272 29850 292300 30049
rect 291200 29786 291252 29792
rect 291304 29804 291382 29832
rect 292260 29844 292312 29850
rect 291212 12034 291240 29786
rect 291200 12028 291252 12034
rect 291200 11970 291252 11976
rect 291304 11966 291332 29804
rect 293173 29832 293201 30049
rect 294091 29832 294119 30049
rect 294992 29832 295020 30049
rect 295910 29832 295938 30049
rect 296794 29866 296822 30049
rect 297712 29866 297740 30049
rect 298647 29866 298675 30049
rect 296794 29838 296852 29866
rect 292260 29786 292312 29792
rect 292592 29804 293201 29832
rect 293972 29804 294119 29832
rect 294984 29804 295020 29832
rect 295904 29804 295938 29832
rect 291844 27396 291896 27402
rect 291844 27338 291896 27344
rect 291856 11966 291884 27338
rect 292592 12102 292620 29804
rect 292580 12096 292632 12102
rect 292580 12038 292632 12044
rect 291292 11960 291344 11966
rect 291292 11902 291344 11908
rect 291844 11960 291896 11966
rect 291844 11902 291896 11908
rect 289820 11892 289872 11898
rect 289820 11834 289872 11840
rect 293972 10878 294000 29804
rect 294984 26234 295012 29804
rect 295904 26234 295932 29804
rect 296076 27328 296128 27334
rect 296076 27270 296128 27276
rect 295984 26308 296036 26314
rect 295984 26250 296036 26256
rect 294064 26206 295012 26234
rect 295352 26206 295932 26234
rect 294064 12170 294092 26206
rect 294604 15020 294656 15026
rect 294604 14962 294656 14968
rect 294052 12164 294104 12170
rect 294052 12106 294104 12112
rect 294512 11892 294564 11898
rect 294512 11834 294564 11840
rect 293960 10872 294012 10878
rect 293960 10814 294012 10820
rect 291384 9444 291436 9450
rect 291384 9386 291436 9392
rect 287060 7948 287112 7954
rect 287060 7890 287112 7896
rect 286600 6452 286652 6458
rect 286600 6394 286652 6400
rect 285680 5296 285732 5302
rect 285680 5238 285732 5244
rect 286612 480 286640 6394
rect 288992 6384 289044 6390
rect 288992 6326 289044 6332
rect 290188 6384 290240 6390
rect 290188 6326 290240 6332
rect 287796 3868 287848 3874
rect 287796 3810 287848 3816
rect 287808 480 287836 3810
rect 289004 480 289032 6326
rect 290200 480 290228 6326
rect 291396 480 291424 9386
rect 292580 6316 292632 6322
rect 292580 6258 292632 6264
rect 293684 6316 293736 6322
rect 293684 6258 293736 6264
rect 292592 480 292620 6258
rect 293696 480 293724 6258
rect 294524 3482 294552 11834
rect 294616 3874 294644 14962
rect 295352 12238 295380 26206
rect 295340 12232 295392 12238
rect 295340 12174 295392 12180
rect 295996 5370 296024 26250
rect 296088 12034 296116 27270
rect 296824 26382 296852 29838
rect 297652 29838 297740 29866
rect 298112 29838 298675 29866
rect 299531 29866 299559 30049
rect 300449 29866 300477 30049
rect 301350 29866 301378 30049
rect 299531 29838 299612 29866
rect 296812 26376 296864 26382
rect 296812 26318 296864 26324
rect 297652 26234 297680 29838
rect 296824 26206 297680 26234
rect 296076 12028 296128 12034
rect 296076 11970 296128 11976
rect 296824 8226 296852 26206
rect 298112 12306 298140 29838
rect 298744 27532 298796 27538
rect 298744 27474 298796 27480
rect 298100 12300 298152 12306
rect 298100 12242 298152 12248
rect 298756 9518 298784 27474
rect 299584 26234 299612 29838
rect 300412 29838 300477 29866
rect 301332 29838 301378 29866
rect 302251 29866 302279 30049
rect 303169 29866 303197 30049
rect 304070 29866 304098 30049
rect 302251 29838 302372 29866
rect 303169 29838 303200 29866
rect 300124 27600 300176 27606
rect 300124 27542 300176 27548
rect 299584 26206 299704 26234
rect 299572 12096 299624 12102
rect 299572 12038 299624 12044
rect 298744 9512 298796 9518
rect 298744 9454 298796 9460
rect 296812 8220 296864 8226
rect 296812 8162 296864 8168
rect 297272 7812 297324 7818
rect 297272 7754 297324 7760
rect 296076 6248 296128 6254
rect 296076 6190 296128 6196
rect 295984 5364 296036 5370
rect 295984 5306 296036 5312
rect 294604 3868 294656 3874
rect 294604 3810 294656 3816
rect 294524 3454 294920 3482
rect 294892 480 294920 3454
rect 296088 480 296116 6190
rect 297284 480 297312 7754
rect 299584 3398 299612 12038
rect 299676 10946 299704 26206
rect 299664 10940 299716 10946
rect 299664 10882 299716 10888
rect 300136 8294 300164 27542
rect 300412 27538 300440 29838
rect 301332 27606 301360 29838
rect 302240 28144 302292 28150
rect 302240 28086 302292 28092
rect 301320 27600 301372 27606
rect 301320 27542 301372 27548
rect 300400 27532 300452 27538
rect 300400 27474 300452 27480
rect 302252 11014 302280 28086
rect 302344 12374 302372 29838
rect 303172 28150 303200 29838
rect 304000 29838 304098 29866
rect 305005 29866 305033 30049
rect 305906 29866 305934 30049
rect 306824 29866 306852 30049
rect 307725 29866 307753 30049
rect 308660 29866 308688 30049
rect 309527 29866 309555 30049
rect 310462 29866 310490 30049
rect 311346 29866 311374 30049
rect 312281 29866 312309 30049
rect 305005 29838 305040 29866
rect 303160 28144 303212 28150
rect 303160 28086 303212 28092
rect 304000 26234 304028 29838
rect 303632 26206 304028 26234
rect 303632 13734 303660 26206
rect 304264 19100 304316 19106
rect 304264 19042 304316 19048
rect 303620 13728 303672 13734
rect 303620 13670 303672 13676
rect 302332 12368 302384 12374
rect 302332 12310 302384 12316
rect 302240 11008 302292 11014
rect 302240 10950 302292 10956
rect 301504 10600 301556 10606
rect 301504 10542 301556 10548
rect 300124 8288 300176 8294
rect 300124 8230 300176 8236
rect 299664 6180 299716 6186
rect 299664 6122 299716 6128
rect 299572 3392 299624 3398
rect 299572 3334 299624 3340
rect 298468 2916 298520 2922
rect 298468 2858 298520 2864
rect 298480 480 298508 2858
rect 299676 480 299704 6122
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300780 480 300808 3334
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 10542
rect 303160 8084 303212 8090
rect 303160 8026 303212 8032
rect 303172 480 303200 8026
rect 304276 2922 304304 19042
rect 305012 6594 305040 29838
rect 305840 29838 305934 29866
rect 306484 29838 306852 29866
rect 307404 29838 307753 29866
rect 308600 29838 308688 29866
rect 309152 29838 309555 29866
rect 310440 29838 310490 29866
rect 311268 29838 311374 29866
rect 311900 29844 311952 29850
rect 305840 26234 305868 29838
rect 306484 26234 306512 29838
rect 307404 26234 307432 29838
rect 308600 26234 308628 29838
rect 305104 26206 305868 26234
rect 306392 26206 306512 26234
rect 306576 26206 307432 26234
rect 307772 26206 308628 26234
rect 305104 6662 305132 26206
rect 306392 6866 306420 26206
rect 306472 23316 306524 23322
rect 306472 23258 306524 23264
rect 306380 6860 306432 6866
rect 306380 6802 306432 6808
rect 305184 6792 305236 6798
rect 305184 6734 305236 6740
rect 305092 6656 305144 6662
rect 305092 6598 305144 6604
rect 305000 6588 305052 6594
rect 305000 6530 305052 6536
rect 304356 6180 304408 6186
rect 304356 6122 304408 6128
rect 304264 2916 304316 2922
rect 304264 2858 304316 2864
rect 304368 480 304396 6122
rect 305196 3806 305224 6734
rect 305552 3936 305604 3942
rect 305552 3878 305604 3884
rect 305184 3800 305236 3806
rect 305184 3742 305236 3748
rect 305564 480 305592 3878
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306484 354 306512 23258
rect 306576 10470 306604 26206
rect 306564 10464 306616 10470
rect 306564 10406 306616 10412
rect 307772 6458 307800 26206
rect 307760 6452 307812 6458
rect 307760 6394 307812 6400
rect 309152 6390 309180 29838
rect 310440 28150 310468 29838
rect 309232 28144 309284 28150
rect 309232 28086 309284 28092
rect 310428 28144 310480 28150
rect 310428 28086 310480 28092
rect 309140 6384 309192 6390
rect 309140 6326 309192 6332
rect 309244 6322 309272 28086
rect 311268 26234 311296 29838
rect 311900 29786 311952 29792
rect 312004 29838 312309 29866
rect 313165 29850 313193 30049
rect 314083 29866 314111 30049
rect 314984 29866 315012 30049
rect 313153 29844 313205 29850
rect 310532 26206 311296 26234
rect 309324 21956 309376 21962
rect 309324 21898 309376 21904
rect 309336 16574 309364 21898
rect 309336 16546 309824 16574
rect 309232 6316 309284 6322
rect 309232 6258 309284 6264
rect 307944 5568 307996 5574
rect 307944 5510 307996 5516
rect 307956 480 307984 5510
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 309060 480 309088 3810
rect 306718 354 306830 480
rect 306484 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 310532 7818 310560 26206
rect 311440 11008 311492 11014
rect 311440 10950 311492 10956
rect 310520 7812 310572 7818
rect 310520 7754 310572 7760
rect 311452 480 311480 10950
rect 311912 6186 311940 29786
rect 312004 12102 312032 29838
rect 313153 29786 313205 29792
rect 313384 29838 314111 29866
rect 314752 29844 314804 29850
rect 312544 25968 312596 25974
rect 312544 25910 312596 25916
rect 311992 12096 312044 12102
rect 311992 12038 312044 12044
rect 311900 6180 311952 6186
rect 311900 6122 311952 6128
rect 312556 3942 312584 25910
rect 313280 24608 313332 24614
rect 313280 24550 313332 24556
rect 312544 3936 312596 3942
rect 312544 3878 312596 3884
rect 312636 3800 312688 3806
rect 312636 3742 312688 3748
rect 312648 480 312676 3742
rect 313292 3482 313320 24550
rect 313384 5574 313412 29838
rect 314752 29786 314804 29792
rect 314948 29838 315012 29866
rect 315902 29850 315930 30049
rect 315890 29844 315942 29850
rect 313924 27600 313976 27606
rect 313924 27542 313976 27548
rect 313936 11014 313964 27542
rect 313924 11008 313976 11014
rect 313924 10950 313976 10956
rect 313372 5568 313424 5574
rect 313372 5510 313424 5516
rect 313292 3454 313872 3482
rect 313844 480 313872 3454
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314764 354 314792 29786
rect 314948 27606 314976 29838
rect 316820 29832 316848 30049
rect 315890 29786 315942 29792
rect 316788 29804 316848 29832
rect 317420 29844 317472 29850
rect 314936 27600 314988 27606
rect 314936 27542 314988 27548
rect 316788 26234 316816 29804
rect 317738 29832 317766 30049
rect 318639 29850 318667 30049
rect 317420 29786 317472 29792
rect 317708 29804 317766 29832
rect 318627 29844 318679 29850
rect 316052 26206 316816 26234
rect 316052 3126 316080 26206
rect 316132 26036 316184 26042
rect 316132 25978 316184 25984
rect 316144 3398 316172 25978
rect 317432 5642 317460 29786
rect 317708 26234 317736 29804
rect 319557 29832 319585 30049
rect 320475 29832 320503 30049
rect 321359 29832 321387 30049
rect 322277 29832 322305 30049
rect 323178 29832 323206 30049
rect 324096 29832 324124 30049
rect 324997 29832 325025 30049
rect 325898 29866 325926 30049
rect 318627 29786 318679 29792
rect 318812 29804 319585 29832
rect 320192 29804 320503 29832
rect 321296 29804 321387 29832
rect 321572 29804 322305 29832
rect 322952 29804 323206 29832
rect 324056 29804 324124 29832
rect 324332 29804 325025 29832
rect 325896 29838 325926 29866
rect 317524 26206 317736 26234
rect 317420 5636 317472 5642
rect 317420 5578 317472 5584
rect 317524 5574 317552 26206
rect 318812 6866 318840 29804
rect 318800 6860 318852 6866
rect 318800 6802 318852 6808
rect 320192 6662 320220 29804
rect 321296 26234 321324 29804
rect 320284 26206 321324 26234
rect 320180 6656 320232 6662
rect 320180 6598 320232 6604
rect 320284 6594 320312 26206
rect 320916 7744 320968 7750
rect 320916 7686 320968 7692
rect 320272 6588 320324 6594
rect 320272 6530 320324 6536
rect 317512 5568 317564 5574
rect 317512 5510 317564 5516
rect 317328 5296 317380 5302
rect 317328 5238 317380 5244
rect 317340 3874 317368 5238
rect 319720 3936 319772 3942
rect 319720 3878 319772 3884
rect 317328 3868 317380 3874
rect 317328 3810 317380 3816
rect 316132 3392 316184 3398
rect 316132 3334 316184 3340
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 316040 3120 316092 3126
rect 316040 3062 316092 3068
rect 316224 3052 316276 3058
rect 316224 2994 316276 3000
rect 316236 480 316264 2994
rect 317340 480 317368 3334
rect 318524 3120 318576 3126
rect 318524 3062 318576 3068
rect 318536 480 318564 3062
rect 319732 480 319760 3878
rect 320928 480 320956 7686
rect 321572 6526 321600 29804
rect 322204 21888 322256 21894
rect 322204 21830 322256 21836
rect 321560 6520 321612 6526
rect 321560 6462 321612 6468
rect 322112 5568 322164 5574
rect 322112 5510 322164 5516
rect 322124 480 322152 5510
rect 322216 3806 322244 21830
rect 322952 6458 322980 29804
rect 324056 26234 324084 29804
rect 323044 26206 324084 26234
rect 322940 6452 322992 6458
rect 322940 6394 322992 6400
rect 323044 6390 323072 26206
rect 323032 6384 323084 6390
rect 323032 6326 323084 6332
rect 324332 6322 324360 29804
rect 325896 27606 325924 29838
rect 325884 27600 325936 27606
rect 325884 27542 325936 27548
rect 326816 26234 326844 30049
rect 327734 29866 327762 30049
rect 328652 29866 328680 30049
rect 329553 29866 329581 30049
rect 330471 29866 330499 30049
rect 331355 29866 331383 30049
rect 332307 29866 332335 30049
rect 333174 29866 333202 30049
rect 334109 29866 334137 30049
rect 334993 29866 335021 30049
rect 335928 29866 335956 30049
rect 327644 29838 327762 29866
rect 328472 29838 328680 29866
rect 328748 29838 329581 29866
rect 329852 29838 330499 29866
rect 331232 29838 331383 29866
rect 331416 29838 332335 29866
rect 333164 29838 333202 29866
rect 333992 29838 334137 29866
rect 334176 29838 335021 29866
rect 335924 29838 335956 29866
rect 336812 29866 336840 30049
rect 337730 29866 337758 30049
rect 338631 29866 338659 30049
rect 336812 29838 336872 29866
rect 327644 26234 327672 29838
rect 327724 27600 327776 27606
rect 327724 27542 327776 27548
rect 325804 26206 326844 26234
rect 327092 26206 327672 26234
rect 325700 20528 325752 20534
rect 325700 20470 325752 20476
rect 324412 17740 324464 17746
rect 324412 17682 324464 17688
rect 324964 17740 325016 17746
rect 324964 17682 325016 17688
rect 324320 6316 324372 6322
rect 324320 6258 324372 6264
rect 322204 3800 322256 3806
rect 322204 3742 322256 3748
rect 323308 3800 323360 3806
rect 323308 3742 323360 3748
rect 323320 480 323348 3742
rect 324424 480 324452 17682
rect 324976 3058 325004 17682
rect 325712 6914 325740 20470
rect 325804 12374 325832 26206
rect 325792 12368 325844 12374
rect 325792 12310 325844 12316
rect 325712 6886 326384 6914
rect 325608 5636 325660 5642
rect 325608 5578 325660 5584
rect 324964 3052 325016 3058
rect 324964 2994 325016 3000
rect 325620 480 325648 5578
rect 314998 354 315110 480
rect 314764 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 6886
rect 327092 6254 327120 26206
rect 327736 12442 327764 27542
rect 327724 12436 327776 12442
rect 327724 12378 327776 12384
rect 328000 12028 328052 12034
rect 328000 11970 328052 11976
rect 327080 6248 327132 6254
rect 327080 6190 327132 6196
rect 328012 480 328040 11970
rect 328472 6186 328500 29838
rect 328748 26234 328776 29838
rect 328564 26206 328776 26234
rect 328564 7954 328592 26206
rect 328552 7948 328604 7954
rect 328552 7890 328604 7896
rect 329852 7886 329880 29838
rect 330484 24608 330536 24614
rect 330484 24550 330536 24556
rect 329840 7880 329892 7886
rect 329840 7822 329892 7828
rect 329196 6860 329248 6866
rect 329196 6802 329248 6808
rect 328460 6180 328512 6186
rect 328460 6122 328512 6128
rect 329208 480 329236 6802
rect 330496 3942 330524 24550
rect 331232 7818 331260 29838
rect 331416 26234 331444 29838
rect 333164 26234 333192 29838
rect 331324 26206 331444 26234
rect 332612 26206 333192 26234
rect 331220 7812 331272 7818
rect 331220 7754 331272 7760
rect 331324 7750 331352 26206
rect 331404 20460 331456 20466
rect 331404 20402 331456 20408
rect 331312 7744 331364 7750
rect 331312 7686 331364 7692
rect 330484 3936 330536 3942
rect 330484 3878 330536 3884
rect 330392 3868 330444 3874
rect 330392 3810 330444 3816
rect 330404 480 330432 3810
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331416 354 331444 20402
rect 332612 8294 332640 26206
rect 332600 8288 332652 8294
rect 332600 8230 332652 8236
rect 333992 8226 334020 29838
rect 334176 26234 334204 29838
rect 335924 26234 335952 29838
rect 336844 27402 336872 29838
rect 337672 29838 337758 29866
rect 338224 29838 338659 29866
rect 339566 29866 339594 30049
rect 340467 29866 340495 30049
rect 341385 29866 341413 30049
rect 342286 29866 342314 30049
rect 343187 29866 343215 30049
rect 344122 29866 344150 30049
rect 339566 29838 339632 29866
rect 336832 27396 336884 27402
rect 336832 27338 336884 27344
rect 337672 26234 337700 29838
rect 334084 26206 334204 26234
rect 335372 26206 335952 26234
rect 336752 26206 337700 26234
rect 334084 11014 334112 26206
rect 334164 19032 334216 19038
rect 334164 18974 334216 18980
rect 334176 16574 334204 18974
rect 334176 16546 334664 16574
rect 334072 11008 334124 11014
rect 334072 10950 334124 10956
rect 333980 8220 334032 8226
rect 333980 8162 334032 8168
rect 332692 6656 332744 6662
rect 332692 6598 332744 6604
rect 332704 480 332732 6598
rect 333888 4004 333940 4010
rect 333888 3946 333940 3952
rect 333900 480 333928 3946
rect 331558 354 331670 480
rect 331416 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335372 10946 335400 26206
rect 336752 23390 336780 26206
rect 338120 24472 338172 24478
rect 338120 24414 338172 24420
rect 336740 23384 336792 23390
rect 336740 23326 336792 23332
rect 336004 15088 336056 15094
rect 336004 15030 336056 15036
rect 335360 10940 335412 10946
rect 335360 10882 335412 10888
rect 336016 3806 336044 15030
rect 338132 6914 338160 24414
rect 338224 10810 338252 29838
rect 339500 28144 339552 28150
rect 339500 28086 339552 28092
rect 339132 27260 339184 27266
rect 339132 27202 339184 27208
rect 339144 24682 339172 27202
rect 339132 24676 339184 24682
rect 339132 24618 339184 24624
rect 338212 10804 338264 10810
rect 338212 10746 338264 10752
rect 339512 10674 339540 28086
rect 339604 10742 339632 29838
rect 340432 29838 340495 29866
rect 341352 29838 341413 29866
rect 342272 29838 342314 29866
rect 342364 29838 343215 29866
rect 344112 29838 344150 29866
rect 345006 29866 345034 30049
rect 345924 29866 345952 30049
rect 346842 29866 346870 30049
rect 345006 29838 345060 29866
rect 340432 28150 340460 29838
rect 340420 28144 340472 28150
rect 340420 28086 340472 28092
rect 341352 27266 341380 29838
rect 341340 27260 341392 27266
rect 341340 27202 341392 27208
rect 341524 23316 341576 23322
rect 341524 23258 341576 23264
rect 340880 23248 340932 23254
rect 340880 23190 340932 23196
rect 339592 10736 339644 10742
rect 339592 10678 339644 10684
rect 339500 10668 339552 10674
rect 339500 10610 339552 10616
rect 338132 6886 338712 6914
rect 337476 6860 337528 6866
rect 337476 6802 337528 6808
rect 336280 6588 336332 6594
rect 336280 6530 336332 6536
rect 336004 3800 336056 3806
rect 336004 3742 336056 3748
rect 336292 480 336320 6530
rect 337488 480 337516 6802
rect 338684 480 338712 6886
rect 339868 6520 339920 6526
rect 339868 6462 339920 6468
rect 339880 480 339908 6462
rect 340892 3398 340920 23190
rect 340972 3936 341024 3942
rect 340972 3878 341024 3884
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 340984 480 341012 3878
rect 341536 3874 341564 23258
rect 342272 19242 342300 29838
rect 342364 21962 342392 29838
rect 344112 26234 344140 29838
rect 343652 26206 344140 26234
rect 343652 26042 343680 26206
rect 343640 26036 343692 26042
rect 343640 25978 343692 25984
rect 342352 21956 342404 21962
rect 342352 21898 342404 21904
rect 342260 19236 342312 19242
rect 342260 19178 342312 19184
rect 345032 17814 345060 29838
rect 345860 29838 345952 29866
rect 346400 29844 346452 29850
rect 345860 26234 345888 29838
rect 346400 29786 346452 29792
rect 346780 29838 346870 29866
rect 347743 29850 347771 30049
rect 348644 29866 348672 30049
rect 349545 29866 349573 30049
rect 350463 29866 350491 30049
rect 351381 29866 351409 30049
rect 352299 29866 352327 30049
rect 347731 29844 347783 29850
rect 345124 26206 345888 26234
rect 345124 24750 345152 26206
rect 345112 24744 345164 24750
rect 345112 24686 345164 24692
rect 345020 17808 345072 17814
rect 345020 17750 345072 17756
rect 342904 16516 342956 16522
rect 342904 16458 342956 16464
rect 342916 4010 342944 16458
rect 346412 13734 346440 29786
rect 346780 26234 346808 29838
rect 347731 29786 347783 29792
rect 348620 29838 348672 29866
rect 349264 29838 349573 29866
rect 349632 29838 350491 29866
rect 350552 29838 351409 29866
rect 352012 29844 352064 29850
rect 348620 27334 348648 29838
rect 348608 27328 348660 27334
rect 348608 27270 348660 27276
rect 346504 26206 346808 26234
rect 346504 20466 346532 26206
rect 349160 21684 349212 21690
rect 349160 21626 349212 21632
rect 346492 20460 346544 20466
rect 346492 20402 346544 20408
rect 346400 13728 346452 13734
rect 346400 13670 346452 13676
rect 345296 11960 345348 11966
rect 345296 11902 345348 11908
rect 343364 6452 343416 6458
rect 343364 6394 343416 6400
rect 342904 4004 342956 4010
rect 342904 3946 342956 3952
rect 341524 3868 341576 3874
rect 341524 3810 341576 3816
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 343376 480 343404 6394
rect 344560 3868 344612 3874
rect 344560 3810 344612 3816
rect 344572 480 344600 3810
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 11902
rect 349172 6914 349200 21626
rect 349264 12306 349292 29838
rect 349632 26234 349660 29838
rect 349356 26206 349660 26234
rect 349252 12300 349304 12306
rect 349252 12242 349304 12248
rect 349356 12238 349384 26206
rect 349344 12232 349396 12238
rect 349344 12174 349396 12180
rect 350552 12170 350580 29838
rect 352012 29786 352064 29792
rect 352116 29838 352327 29866
rect 353200 29850 353228 30049
rect 354135 29866 354163 30049
rect 355002 29866 355030 30049
rect 353188 29844 353240 29850
rect 351920 25900 351972 25906
rect 351920 25842 351972 25848
rect 350540 12164 350592 12170
rect 350540 12106 350592 12112
rect 351932 6914 351960 25842
rect 352024 12034 352052 29786
rect 352116 12102 352144 29838
rect 353188 29786 353240 29792
rect 353312 29838 354163 29866
rect 354968 29838 355030 29866
rect 355954 29866 355982 30049
rect 356821 29866 356849 30049
rect 357756 29866 357784 30049
rect 355954 29838 356008 29866
rect 352104 12096 352156 12102
rect 352104 12038 352156 12044
rect 352012 12028 352064 12034
rect 352012 11970 352064 11976
rect 353312 11966 353340 29838
rect 353392 27396 353444 27402
rect 353392 27338 353444 27344
rect 353404 26178 353432 27338
rect 354968 26234 354996 29838
rect 355980 27606 356008 29838
rect 356072 29838 356849 29866
rect 357440 29844 357492 29850
rect 355968 27600 356020 27606
rect 355968 27542 356020 27548
rect 354692 26206 354996 26234
rect 353392 26172 353444 26178
rect 353392 26114 353444 26120
rect 354692 23254 354720 26206
rect 356072 25906 356100 29838
rect 357440 29786 357492 29792
rect 357728 29838 357784 29866
rect 358657 29850 358685 30049
rect 359575 29866 359603 30049
rect 360459 29866 360487 30049
rect 358645 29844 358697 29850
rect 356704 27600 356756 27606
rect 356704 27542 356756 27548
rect 356060 25900 356112 25906
rect 356060 25842 356112 25848
rect 354680 23248 354732 23254
rect 354680 23190 354732 23196
rect 353944 19032 353996 19038
rect 353944 18974 353996 18980
rect 353576 12436 353628 12442
rect 353576 12378 353628 12384
rect 353300 11960 353352 11966
rect 353300 11902 353352 11908
rect 349172 6886 349292 6914
rect 351932 6886 352880 6914
rect 346952 6384 347004 6390
rect 346952 6326 347004 6332
rect 346964 480 346992 6326
rect 348056 5364 348108 5370
rect 348056 5306 348108 5312
rect 348068 480 348096 5306
rect 349264 480 349292 6886
rect 350448 6316 350500 6322
rect 350448 6258 350500 6264
rect 350460 480 350488 6258
rect 351644 3800 351696 3806
rect 351644 3742 351696 3748
rect 351656 480 351684 3742
rect 352852 480 352880 6886
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 12378
rect 353956 3942 353984 18974
rect 356716 9518 356744 27542
rect 356704 9512 356756 9518
rect 356704 9454 356756 9460
rect 356336 7676 356388 7682
rect 356336 7618 356388 7624
rect 356060 7540 356112 7546
rect 356060 7482 356112 7488
rect 355232 4004 355284 4010
rect 355232 3946 355284 3952
rect 353944 3936 353996 3942
rect 353944 3878 353996 3884
rect 355244 480 355272 3946
rect 356072 3738 356100 7482
rect 356060 3732 356112 3738
rect 356060 3674 356112 3680
rect 356348 480 356376 7618
rect 357452 6662 357480 29786
rect 357728 26234 357756 29838
rect 358645 29786 358697 29792
rect 358832 29838 359603 29866
rect 360212 29838 360487 29866
rect 361377 29866 361405 30049
rect 362278 29866 362306 30049
rect 363213 29866 363241 30049
rect 361377 29838 361436 29866
rect 362278 29838 362356 29866
rect 357544 26206 357756 26234
rect 357544 16454 357572 26206
rect 357532 16448 357584 16454
rect 357532 16390 357584 16396
rect 357532 12368 357584 12374
rect 357532 12310 357584 12316
rect 357440 6656 357492 6662
rect 357440 6598 357492 6604
rect 357544 480 357572 12310
rect 358832 6594 358860 29838
rect 358912 17672 358964 17678
rect 358912 17614 358964 17620
rect 358924 16574 358952 17614
rect 358924 16546 359504 16574
rect 358820 6588 358872 6594
rect 358820 6530 358872 6536
rect 358728 3732 358780 3738
rect 358728 3674 358780 3680
rect 358740 480 358768 3674
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 360212 6526 360240 29838
rect 361408 27538 361436 29838
rect 361396 27532 361448 27538
rect 361396 27474 361448 27480
rect 362328 27402 362356 29838
rect 362960 29844 363012 29850
rect 362960 29786 363012 29792
rect 363064 29838 363241 29866
rect 364114 29850 364142 30049
rect 365032 29866 365060 30049
rect 364102 29844 364154 29850
rect 362316 27396 362368 27402
rect 362316 27338 362368 27344
rect 360476 27260 360528 27266
rect 360476 27202 360528 27208
rect 360488 20602 360516 27202
rect 360476 20596 360528 20602
rect 360476 20538 360528 20544
rect 360844 13048 360896 13054
rect 360844 12990 360896 12996
rect 360200 6520 360252 6526
rect 360200 6462 360252 6468
rect 360856 3874 360884 12990
rect 362972 6390 363000 29786
rect 363064 6458 363092 29838
rect 364102 29786 364154 29792
rect 364904 29838 365060 29866
rect 364904 26234 364932 29838
rect 365950 29832 365978 30049
rect 366834 29832 366862 30049
rect 367769 29832 367797 30049
rect 365732 29804 365978 29832
rect 366744 29804 366862 29832
rect 367112 29804 367797 29832
rect 364984 27328 365036 27334
rect 364984 27270 365036 27276
rect 364352 26206 364932 26234
rect 363144 20324 363196 20330
rect 363144 20266 363196 20272
rect 363156 16574 363184 20266
rect 363156 16546 363552 16574
rect 363052 6452 363104 6458
rect 363052 6394 363104 6400
rect 362960 6384 363012 6390
rect 362960 6326 363012 6332
rect 361120 6248 361172 6254
rect 361120 6190 361172 6196
rect 360844 3868 360896 3874
rect 360844 3810 360896 3816
rect 361132 480 361160 6190
rect 362316 4072 362368 4078
rect 362316 4014 362368 4020
rect 362328 480 362356 4014
rect 363524 480 363552 16546
rect 364352 6322 364380 26206
rect 364996 19174 365024 27270
rect 364984 19168 365036 19174
rect 364984 19110 365036 19116
rect 364340 6316 364392 6322
rect 364340 6258 364392 6264
rect 365732 6254 365760 29804
rect 366744 26234 366772 29804
rect 365824 26206 366772 26234
rect 365720 6248 365772 6254
rect 365720 6190 365772 6196
rect 365824 6186 365852 26206
rect 367112 24478 367140 29804
rect 368653 29730 368681 30049
rect 369571 29832 369599 30049
rect 370489 29832 370517 30049
rect 371390 29832 371418 30049
rect 372291 29832 372319 30049
rect 373209 29832 373237 30049
rect 374110 29866 374138 30049
rect 368768 29804 369599 29832
rect 369964 29804 370517 29832
rect 371252 29804 371418 29832
rect 371620 29804 372319 29832
rect 372632 29804 373237 29832
rect 374000 29844 374052 29850
rect 368653 29702 368704 29730
rect 368676 27470 368704 29702
rect 368664 27464 368716 27470
rect 368664 27406 368716 27412
rect 367744 27328 367796 27334
rect 367744 27270 367796 27276
rect 367100 24472 367152 24478
rect 367100 24414 367152 24420
rect 365904 18964 365956 18970
rect 365904 18906 365956 18912
rect 365916 16574 365944 18906
rect 365916 16546 367048 16574
rect 364616 6180 364668 6186
rect 364616 6122 364668 6128
rect 365812 6180 365864 6186
rect 365812 6122 365864 6128
rect 364628 480 364656 6122
rect 365812 3868 365864 3874
rect 365812 3810 365864 3816
rect 365824 480 365852 3810
rect 367020 480 367048 16546
rect 367756 6730 367784 27270
rect 368768 26234 368796 29804
rect 368492 26206 368796 26234
rect 367836 22024 367888 22030
rect 367836 21966 367888 21972
rect 367744 6724 367796 6730
rect 367744 6666 367796 6672
rect 367848 3806 367876 21966
rect 368492 9382 368520 26206
rect 369860 24404 369912 24410
rect 369860 24346 369912 24352
rect 368480 9376 368532 9382
rect 368480 9318 368532 9324
rect 368204 7948 368256 7954
rect 368204 7890 368256 7896
rect 367836 3800 367888 3806
rect 367836 3742 367888 3748
rect 368216 480 368244 7890
rect 369872 6914 369900 24346
rect 369964 13462 369992 29804
rect 369952 13456 370004 13462
rect 369952 13398 370004 13404
rect 371252 10470 371280 29804
rect 371620 26234 371648 29804
rect 371344 26206 371648 26234
rect 371344 23050 371372 26206
rect 371332 23044 371384 23050
rect 371332 22986 371384 22992
rect 372632 21690 372660 29804
rect 374000 29786 374052 29792
rect 374104 29838 374138 29866
rect 375028 29850 375056 30049
rect 375946 29866 375974 30049
rect 375016 29844 375068 29850
rect 372620 21684 372672 21690
rect 372620 21626 372672 21632
rect 374012 16114 374040 29786
rect 374104 17678 374132 29838
rect 375016 29786 375068 29792
rect 375944 29838 375974 29866
rect 376847 29866 376875 30049
rect 377782 29866 377810 30049
rect 378649 29866 378677 30049
rect 376847 29838 376892 29866
rect 375944 26234 375972 29838
rect 376116 27532 376168 27538
rect 376116 27474 376168 27480
rect 375392 26206 375972 26234
rect 374092 17672 374144 17678
rect 374092 17614 374144 17620
rect 374000 16108 374052 16114
rect 374000 16050 374052 16056
rect 374092 13660 374144 13666
rect 374092 13602 374144 13608
rect 371240 10464 371292 10470
rect 371240 10406 371292 10412
rect 371700 7880 371752 7886
rect 371700 7822 371752 7828
rect 369872 6886 370176 6914
rect 369400 3800 369452 3806
rect 369400 3742 369452 3748
rect 369412 480 369440 3742
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 354 370176 6886
rect 371712 480 371740 7822
rect 372896 3936 372948 3942
rect 372896 3878 372948 3884
rect 372908 480 372936 3878
rect 374104 480 374132 13602
rect 375392 8090 375420 26206
rect 376024 26104 376076 26110
rect 376024 26046 376076 26052
rect 375380 8084 375432 8090
rect 375380 8026 375432 8032
rect 375288 7812 375340 7818
rect 375288 7754 375340 7760
rect 375300 480 375328 7754
rect 376036 4010 376064 26046
rect 376128 13598 376156 27474
rect 376760 23112 376812 23118
rect 376760 23054 376812 23060
rect 376116 13592 376168 13598
rect 376116 13534 376168 13540
rect 376772 6914 376800 23054
rect 376864 8022 376892 29838
rect 377692 29838 377810 29866
rect 378152 29838 378677 29866
rect 377692 26234 377720 29838
rect 376956 26206 377720 26234
rect 376852 8016 376904 8022
rect 376852 7958 376904 7964
rect 376956 7954 376984 26206
rect 376944 7948 376996 7954
rect 376944 7890 376996 7896
rect 378152 7886 378180 29838
rect 379584 29832 379612 30049
rect 380468 29832 380496 30049
rect 381403 29832 381431 30049
rect 379584 29804 379652 29832
rect 379624 26382 379652 29804
rect 380452 29804 380496 29832
rect 380912 29804 381431 29832
rect 382304 29832 382332 30049
rect 383222 29832 383250 30049
rect 384106 29832 384134 30049
rect 382304 29804 382412 29832
rect 380452 27266 380480 29804
rect 380440 27260 380492 27266
rect 380440 27202 380492 27208
rect 379612 26376 379664 26382
rect 379612 26318 379664 26324
rect 378784 15156 378836 15162
rect 378784 15098 378836 15104
rect 378140 7880 378192 7886
rect 378140 7822 378192 7828
rect 376772 6886 377720 6914
rect 376484 4140 376536 4146
rect 376484 4082 376536 4088
rect 376024 4004 376076 4010
rect 376024 3946 376076 3952
rect 376496 480 376524 4082
rect 377692 480 377720 6886
rect 378796 4078 378824 15098
rect 380912 7818 380940 29804
rect 381544 26376 381596 26382
rect 381544 26318 381596 26324
rect 380992 21752 381044 21758
rect 380992 21694 381044 21700
rect 381004 16574 381032 21694
rect 381004 16546 381216 16574
rect 380900 7812 380952 7818
rect 380900 7754 380952 7760
rect 378876 7744 378928 7750
rect 378876 7686 378928 7692
rect 378784 4072 378836 4078
rect 378784 4014 378836 4020
rect 378888 480 378916 7686
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 379992 480 380020 3946
rect 381188 480 381216 16546
rect 381556 14890 381584 26318
rect 382280 26240 382332 26246
rect 382280 26182 382332 26188
rect 381544 14884 381596 14890
rect 381544 14826 381596 14832
rect 381544 10872 381596 10878
rect 381544 10814 381596 10820
rect 381556 3738 381584 10814
rect 382292 7682 382320 26182
rect 382384 16574 382412 29804
rect 383212 29804 383250 29832
rect 384040 29804 384134 29832
rect 385041 29832 385069 30049
rect 385925 29832 385953 30049
rect 386860 29832 386888 30049
rect 387761 29866 387789 30049
rect 385041 29804 385080 29832
rect 383212 26246 383240 29804
rect 383200 26240 383252 26246
rect 383200 26182 383252 26188
rect 383660 25832 383712 25838
rect 383660 25774 383712 25780
rect 382384 16546 382504 16574
rect 382372 8288 382424 8294
rect 382372 8230 382424 8236
rect 382280 7676 382332 7682
rect 382280 7618 382332 7624
rect 381544 3732 381596 3738
rect 381544 3674 381596 3680
rect 382384 480 382412 8230
rect 382476 7750 382504 16546
rect 382464 7744 382516 7750
rect 382464 7686 382516 7692
rect 383672 6914 383700 25774
rect 384040 22094 384068 29804
rect 383764 22066 384068 22094
rect 383764 13122 383792 22066
rect 383752 13116 383804 13122
rect 383752 13058 383804 13064
rect 385052 7614 385080 29804
rect 385144 29804 385953 29832
rect 386800 29804 386888 29832
rect 387720 29838 387789 29866
rect 385144 14482 385172 29804
rect 386420 26240 386472 26246
rect 386420 26182 386472 26188
rect 385684 24404 385736 24410
rect 385684 24346 385736 24352
rect 385132 14476 385184 14482
rect 385132 14418 385184 14424
rect 385040 7608 385092 7614
rect 385040 7550 385092 7556
rect 383672 6886 384344 6914
rect 383566 3360 383622 3369
rect 383566 3295 383622 3304
rect 383580 480 383608 3295
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 6886
rect 385696 4146 385724 24346
rect 385960 8220 386012 8226
rect 385960 8162 386012 8168
rect 385684 4140 385736 4146
rect 385684 4082 385736 4088
rect 385972 480 386000 8162
rect 386432 6798 386460 26182
rect 386800 22094 386828 29804
rect 387720 26246 387748 29838
rect 388679 29832 388707 30049
rect 389597 29866 389625 30049
rect 388272 29804 388707 29832
rect 389180 29844 389232 29850
rect 387708 26240 387760 26246
rect 387708 26182 387760 26188
rect 388272 22094 388300 29804
rect 389180 29786 389232 29792
rect 389284 29838 389625 29866
rect 390481 29850 390509 30049
rect 391399 29866 391427 30049
rect 392317 29866 392345 30049
rect 390469 29844 390521 29850
rect 386524 22066 386828 22094
rect 387812 22066 388300 22094
rect 386524 15910 386552 22066
rect 386512 15904 386564 15910
rect 386512 15846 386564 15852
rect 387812 7546 387840 22066
rect 387892 17604 387944 17610
rect 387892 17546 387944 17552
rect 387800 7540 387852 7546
rect 387800 7482 387852 7488
rect 386420 6792 386472 6798
rect 386420 6734 386472 6740
rect 387156 3732 387208 3738
rect 387156 3674 387208 3680
rect 387168 480 387196 3674
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387904 354 387932 17546
rect 389192 3534 389220 29786
rect 389180 3528 389232 3534
rect 389180 3470 389232 3476
rect 389284 3466 389312 29838
rect 390469 29786 390521 29792
rect 390572 29838 391427 29866
rect 392136 29838 392345 29866
rect 393218 29866 393246 30049
rect 394136 29866 394164 30049
rect 395037 29866 395065 30049
rect 395938 29866 395966 30049
rect 396856 29866 396884 30049
rect 397757 29866 397785 30049
rect 398675 29866 398703 30049
rect 399593 29866 399621 30049
rect 400477 29866 400505 30049
rect 401429 29866 401457 30049
rect 402296 29866 402324 30049
rect 403231 29866 403259 30049
rect 404132 29866 404160 30049
rect 405050 29866 405078 30049
rect 405951 29866 405979 30049
rect 393218 29838 393268 29866
rect 389456 11008 389508 11014
rect 389456 10950 389508 10956
rect 389272 3460 389324 3466
rect 389272 3402 389324 3408
rect 389468 480 389496 10950
rect 390572 3602 390600 29838
rect 390652 24676 390704 24682
rect 390652 24618 390704 24624
rect 390560 3596 390612 3602
rect 390560 3538 390612 3544
rect 390664 3534 390692 24618
rect 392032 10940 392084 10946
rect 392032 10882 392084 10888
rect 390652 3528 390704 3534
rect 390652 3470 390704 3476
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 390664 480 390692 3334
rect 391860 480 391888 3470
rect 392044 490 392072 10882
rect 392136 3670 392164 29838
rect 393240 28286 393268 29838
rect 394068 29838 394164 29866
rect 394712 29838 395065 29866
rect 395908 29838 395966 29866
rect 396828 29838 396884 29866
rect 397748 29838 397785 29866
rect 398668 29838 398703 29866
rect 399036 29838 399621 29866
rect 400416 29838 400505 29866
rect 401428 29838 401457 29866
rect 402256 29838 402324 29866
rect 403176 29838 403259 29866
rect 403544 29838 404160 29866
rect 405016 29838 405078 29866
rect 405740 29844 405792 29850
rect 393228 28280 393280 28286
rect 393228 28222 393280 28228
rect 394068 26234 394096 29838
rect 393332 26206 394096 26234
rect 392124 3664 392176 3670
rect 392124 3606 392176 3612
rect 393332 2174 393360 26206
rect 394712 13190 394740 29838
rect 395908 26234 395936 29838
rect 396828 28354 396856 29838
rect 396816 28348 396868 28354
rect 396816 28290 396868 28296
rect 397748 27606 397776 29838
rect 398668 28422 398696 29838
rect 398656 28416 398708 28422
rect 398656 28358 398708 28364
rect 396724 27600 396776 27606
rect 396724 27542 396776 27548
rect 397736 27600 397788 27606
rect 397736 27542 397788 27548
rect 394804 26206 395936 26234
rect 394804 13258 394832 26206
rect 396080 26172 396132 26178
rect 396080 26114 396132 26120
rect 394884 20256 394936 20262
rect 394884 20198 394936 20204
rect 394896 16574 394924 20198
rect 394896 16546 395384 16574
rect 394792 13252 394844 13258
rect 394792 13194 394844 13200
rect 394700 13184 394752 13190
rect 394700 13126 394752 13132
rect 394240 3392 394292 3398
rect 394240 3334 394292 3340
rect 393320 2168 393372 2174
rect 393320 2110 393372 2116
rect 388230 354 388342 480
rect 387904 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392044 462 392624 490
rect 394252 480 394280 3334
rect 395356 480 395384 16546
rect 392596 354 392624 462
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 26114
rect 396736 2242 396764 27542
rect 396816 27124 396868 27130
rect 396816 27066 396868 27072
rect 396828 13122 396856 27066
rect 398840 23384 398892 23390
rect 398840 23326 398892 23332
rect 396816 13116 396868 13122
rect 396816 13058 396868 13064
rect 397736 3596 397788 3602
rect 397736 3538 397788 3544
rect 396724 2236 396776 2242
rect 396724 2178 396776 2184
rect 397748 480 397776 3538
rect 398852 3534 398880 23326
rect 398932 18896 398984 18902
rect 398932 18838 398984 18844
rect 398840 3528 398892 3534
rect 398840 3470 398892 3476
rect 398944 480 398972 18838
rect 399036 11762 399064 29838
rect 399024 11756 399076 11762
rect 399024 11698 399076 11704
rect 400128 3528 400180 3534
rect 400128 3470 400180 3476
rect 400140 480 400168 3470
rect 400416 2310 400444 29838
rect 401428 28490 401456 29838
rect 401416 28484 401468 28490
rect 401416 28426 401468 28432
rect 402256 26234 402284 29838
rect 403176 28558 403204 29838
rect 403164 28552 403216 28558
rect 403164 28494 403216 28500
rect 403544 26234 403572 29838
rect 403624 27124 403676 27130
rect 403624 27066 403676 27072
rect 401612 26206 402284 26234
rect 403084 26206 403572 26234
rect 400680 9580 400732 9586
rect 400680 9522 400732 9528
rect 400692 3874 400720 9522
rect 400680 3868 400732 3874
rect 400680 3810 400732 3816
rect 401324 3664 401376 3670
rect 401324 3606 401376 3612
rect 400404 2304 400456 2310
rect 400404 2246 400456 2252
rect 401336 480 401364 3606
rect 401612 2378 401640 26206
rect 403084 14550 403112 26206
rect 403072 14544 403124 14550
rect 403072 14486 403124 14492
rect 403532 10804 403584 10810
rect 403532 10746 403584 10752
rect 402520 9308 402572 9314
rect 402520 9250 402572 9256
rect 401600 2372 401652 2378
rect 401600 2314 401652 2320
rect 402532 480 402560 9250
rect 403544 3482 403572 10746
rect 403636 6866 403664 27066
rect 405016 26234 405044 29838
rect 405740 29786 405792 29792
rect 405844 29838 405979 29866
rect 406869 29850 406897 30049
rect 407753 29866 407781 30049
rect 406857 29844 406909 29850
rect 404372 26206 405044 26234
rect 404372 14618 404400 26206
rect 405752 14754 405780 29786
rect 405740 14748 405792 14754
rect 405740 14690 405792 14696
rect 405844 14686 405872 29838
rect 406857 29786 406909 29792
rect 407132 29838 407781 29866
rect 408671 29866 408699 30049
rect 409572 29866 409600 30049
rect 410473 29866 410501 30049
rect 411374 29866 411402 30049
rect 412292 29866 412320 30049
rect 408671 29838 408724 29866
rect 407132 14822 407160 29838
rect 408696 27606 408724 29838
rect 409524 29838 409600 29866
rect 409892 29838 410501 29866
rect 411272 29838 411402 29866
rect 412284 29838 412320 29866
rect 407764 27600 407816 27606
rect 407764 27542 407816 27548
rect 408684 27600 408736 27606
rect 408684 27542 408736 27548
rect 407120 14816 407172 14822
rect 407120 14758 407172 14764
rect 405832 14680 405884 14686
rect 405832 14622 405884 14628
rect 404360 14612 404412 14618
rect 404360 14554 404412 14560
rect 405004 14612 405056 14618
rect 405004 14554 405056 14560
rect 403716 10804 403768 10810
rect 403716 10746 403768 10752
rect 403624 6860 403676 6866
rect 403624 6802 403676 6808
rect 403728 3806 403756 10746
rect 405016 3942 405044 14554
rect 407212 10736 407264 10742
rect 407212 10678 407264 10684
rect 406016 9240 406068 9246
rect 406016 9182 406068 9188
rect 405004 3936 405056 3942
rect 405004 3878 405056 3884
rect 403716 3800 403768 3806
rect 403716 3742 403768 3748
rect 404820 3800 404872 3806
rect 404820 3742 404872 3748
rect 403544 3454 403664 3482
rect 403636 480 403664 3454
rect 404832 480 404860 3742
rect 406028 480 406056 9182
rect 407224 480 407252 10678
rect 407776 5234 407804 27542
rect 407856 27192 407908 27198
rect 407856 27134 407908 27140
rect 407868 14482 407896 27134
rect 409524 26234 409552 29838
rect 408604 26206 409552 26234
rect 408604 17542 408632 26206
rect 408592 17536 408644 17542
rect 408592 17478 408644 17484
rect 409892 14958 409920 29838
rect 410524 27396 410576 27402
rect 410524 27338 410576 27344
rect 410432 27192 410484 27198
rect 410432 27134 410484 27140
rect 410444 21826 410472 27134
rect 410432 21820 410484 21826
rect 410432 21762 410484 21768
rect 409880 14952 409932 14958
rect 409880 14894 409932 14900
rect 410536 14550 410564 27338
rect 410524 14544 410576 14550
rect 410524 14486 410576 14492
rect 407856 14476 407908 14482
rect 407856 14418 407908 14424
rect 410800 10668 410852 10674
rect 410800 10610 410852 10616
rect 409604 9172 409656 9178
rect 409604 9114 409656 9120
rect 407764 5228 407816 5234
rect 407764 5170 407816 5176
rect 408408 3868 408460 3874
rect 408408 3810 408460 3816
rect 408420 480 408448 3810
rect 409616 480 409644 9114
rect 410812 480 410840 10610
rect 411272 10538 411300 29838
rect 412284 26234 412312 29838
rect 413210 29832 413238 30049
rect 414111 29832 414139 30049
rect 415029 29832 415057 30049
rect 413204 29804 413238 29832
rect 414032 29804 414139 29832
rect 414492 29804 415057 29832
rect 415947 29832 415975 30049
rect 416848 29832 416876 30049
rect 417766 29832 417794 30049
rect 418684 29832 418712 30049
rect 415947 29804 415992 29832
rect 413204 26234 413232 29804
rect 413284 27396 413336 27402
rect 413284 27338 413336 27344
rect 411364 26206 412312 26234
rect 412744 26206 413232 26234
rect 411364 15978 411392 26206
rect 412640 24336 412692 24342
rect 412640 24278 412692 24284
rect 411904 16584 411956 16590
rect 411904 16526 411956 16532
rect 411352 15972 411404 15978
rect 411352 15914 411404 15920
rect 411260 10532 411312 10538
rect 411260 10474 411312 10480
rect 411916 4078 411944 16526
rect 411904 4072 411956 4078
rect 411904 4014 411956 4020
rect 411904 3936 411956 3942
rect 411904 3878 411956 3884
rect 411916 480 411944 3878
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 24278
rect 412744 16046 412772 26206
rect 412732 16040 412784 16046
rect 412732 15982 412784 15988
rect 413296 11898 413324 27338
rect 414032 16182 414060 29804
rect 414492 26234 414520 29804
rect 414664 27464 414716 27470
rect 414664 27406 414716 27412
rect 414124 26206 414520 26234
rect 414124 16250 414152 26206
rect 414204 20596 414256 20602
rect 414204 20538 414256 20544
rect 414216 16574 414244 20538
rect 414216 16546 414336 16574
rect 414112 16244 414164 16250
rect 414112 16186 414164 16192
rect 414020 16176 414072 16182
rect 414020 16118 414072 16124
rect 413284 11892 413336 11898
rect 413284 11834 413336 11840
rect 414308 480 414336 16546
rect 414676 15910 414704 27406
rect 415964 27198 415992 29804
rect 416792 29804 416876 29832
rect 417712 29804 417794 29832
rect 418632 29804 418712 29832
rect 419534 29832 419562 30049
rect 420486 29832 420514 30049
rect 421353 29832 421381 30049
rect 419534 29804 419580 29832
rect 416688 27600 416740 27606
rect 416688 27542 416740 27548
rect 415952 27192 416004 27198
rect 415952 27134 416004 27140
rect 416700 23186 416728 27542
rect 416688 23180 416740 23186
rect 416688 23122 416740 23128
rect 416792 16318 416820 29804
rect 417712 26234 417740 29804
rect 418632 26234 418660 29804
rect 419552 27334 419580 29804
rect 420472 29804 420514 29832
rect 421300 29804 421381 29832
rect 422288 29832 422316 30049
rect 423206 29832 423234 30049
rect 424107 29832 424135 30049
rect 422288 29804 422340 29832
rect 419540 27328 419592 27334
rect 419540 27270 419592 27276
rect 418804 27192 418856 27198
rect 418804 27134 418856 27140
rect 416884 26206 417740 26234
rect 418172 26206 418660 26234
rect 416884 16386 416912 26206
rect 416964 19236 417016 19242
rect 416964 19178 417016 19184
rect 416976 16574 417004 19178
rect 416976 16546 417464 16574
rect 416872 16380 416924 16386
rect 416872 16322 416924 16328
rect 416780 16312 416832 16318
rect 416780 16254 416832 16260
rect 414664 15904 414716 15910
rect 414664 15846 414716 15852
rect 415400 13388 415452 13394
rect 415400 13330 415452 13336
rect 415412 3398 415440 13330
rect 415492 4004 415544 4010
rect 415492 3946 415544 3952
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 3946
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418172 11830 418200 26206
rect 418160 11824 418212 11830
rect 418160 11766 418212 11772
rect 418816 5370 418844 27134
rect 418896 27056 418948 27062
rect 418896 26998 418948 27004
rect 418908 15978 418936 26998
rect 420472 26234 420500 29804
rect 421300 27606 421328 29804
rect 421288 27600 421340 27606
rect 421288 27542 421340 27548
rect 421564 27056 421616 27062
rect 421564 26998 421616 27004
rect 421012 26308 421064 26314
rect 421012 26250 421064 26256
rect 419644 26206 420500 26234
rect 419644 24546 419672 26206
rect 419632 24540 419684 24546
rect 419632 24482 419684 24488
rect 420920 21956 420972 21962
rect 420920 21898 420972 21904
rect 418896 15972 418948 15978
rect 418896 15914 418948 15920
rect 420184 9104 420236 9110
rect 420184 9046 420236 9052
rect 418804 5364 418856 5370
rect 418804 5306 418856 5312
rect 418988 4072 419040 4078
rect 418988 4014 419040 4020
rect 419000 480 419028 4014
rect 420196 480 420224 9046
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 21898
rect 421024 20398 421052 26250
rect 421012 20392 421064 20398
rect 421012 20334 421064 20340
rect 421576 9450 421604 26998
rect 421564 9444 421616 9450
rect 421564 9386 421616 9392
rect 422312 8158 422340 29804
rect 423140 29804 423234 29832
rect 424060 29804 424135 29832
rect 425042 29832 425070 30049
rect 425926 29832 425954 30049
rect 425042 29804 425100 29832
rect 423140 26234 423168 29804
rect 424060 26314 424088 29804
rect 424324 26988 424376 26994
rect 424324 26930 424376 26936
rect 424416 26988 424468 26994
rect 424416 26930 424468 26936
rect 424048 26308 424100 26314
rect 424048 26250 424100 26256
rect 422404 26206 423168 26234
rect 422404 13530 422432 26206
rect 423680 26036 423732 26042
rect 423680 25978 423732 25984
rect 422392 13524 422444 13530
rect 422392 13466 422444 13472
rect 422300 8152 422352 8158
rect 422300 8094 422352 8100
rect 422576 4140 422628 4146
rect 422576 4082 422628 4088
rect 422588 480 422616 4082
rect 423692 3398 423720 25978
rect 424336 9042 424364 26930
rect 424428 20534 424456 26930
rect 425072 26234 425100 29804
rect 425900 29804 425954 29832
rect 426532 29844 426584 29850
rect 425704 27600 425756 27606
rect 425704 27542 425756 27548
rect 425072 26206 425192 26234
rect 424416 20528 424468 20534
rect 424416 20470 424468 20476
rect 425164 15026 425192 26206
rect 425152 15020 425204 15026
rect 425152 14962 425204 14968
rect 425716 10606 425744 27542
rect 425900 27062 425928 29804
rect 426861 29832 426889 30049
rect 427762 29850 427790 30049
rect 426532 29786 426584 29792
rect 426820 29804 426889 29832
rect 427750 29844 427802 29850
rect 425888 27056 425940 27062
rect 425888 26998 425940 27004
rect 426440 22976 426492 22982
rect 426440 22918 426492 22924
rect 426452 16574 426480 22918
rect 426544 19106 426572 29786
rect 426820 27402 426848 29804
rect 428680 29832 428708 30049
rect 429581 29832 429609 30049
rect 430516 29832 430544 30049
rect 431366 29832 431394 30049
rect 432318 29866 432346 30049
rect 427750 29786 427802 29792
rect 428660 29804 428708 29832
rect 429212 29804 429609 29832
rect 430500 29804 430544 29832
rect 431328 29804 431394 29832
rect 431960 29844 432012 29850
rect 428660 27606 428688 29804
rect 428648 27600 428700 27606
rect 428648 27542 428700 27548
rect 426808 27396 426860 27402
rect 426808 27338 426860 27344
rect 428464 26920 428516 26926
rect 428464 26862 428516 26868
rect 426532 19100 426584 19106
rect 426532 19042 426584 19048
rect 427820 17808 427872 17814
rect 427820 17750 427872 17756
rect 426452 16546 426848 16574
rect 425704 10600 425756 10606
rect 425704 10542 425756 10548
rect 423772 9036 423824 9042
rect 423772 8978 423824 8984
rect 424324 9036 424376 9042
rect 424324 8978 424376 8984
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 8978
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 426164 3392 426216 3398
rect 426164 3334 426216 3340
rect 424980 480 425008 3334
rect 426176 480 426204 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 427832 6914 427860 17750
rect 428476 8362 428504 26862
rect 429212 25974 429240 29804
rect 430500 28150 430528 29804
rect 429292 28144 429344 28150
rect 429292 28086 429344 28092
rect 430488 28144 430540 28150
rect 430488 28086 430540 28092
rect 429200 25968 429252 25974
rect 429200 25910 429252 25916
rect 428464 8356 428516 8362
rect 428464 8298 428516 8304
rect 427832 6886 428504 6914
rect 428476 480 428504 6886
rect 429304 5302 429332 28086
rect 429384 26920 429436 26926
rect 429384 26862 429436 26868
rect 429292 5296 429344 5302
rect 429292 5238 429344 5244
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429396 354 429424 26862
rect 431328 26234 431356 29804
rect 431960 29786 432012 29792
rect 432248 29838 432346 29866
rect 433185 29850 433213 30049
rect 434120 29866 434148 30049
rect 435021 29866 435049 30049
rect 433173 29844 433225 29850
rect 430592 26206 431356 26234
rect 430592 21894 430620 26206
rect 431972 24614 432000 29786
rect 432248 26234 432276 29838
rect 433173 29786 433225 29792
rect 434088 29838 434148 29866
rect 434812 29844 434864 29850
rect 434088 26234 434116 29838
rect 434812 29786 434864 29792
rect 435008 29838 435049 29866
rect 435939 29850 435967 30049
rect 436857 29866 436885 30049
rect 437775 29866 437803 30049
rect 438676 29866 438704 30049
rect 439594 29866 439622 30049
rect 440495 29866 440523 30049
rect 441413 29866 441441 30049
rect 442331 29866 442359 30049
rect 443181 29866 443209 30049
rect 444133 29866 444161 30049
rect 445034 29866 445062 30049
rect 445935 29866 445963 30049
rect 446853 29866 446881 30049
rect 447754 29866 447782 30049
rect 448689 29866 448717 30049
rect 435927 29844 435979 29850
rect 432064 26206 432276 26234
rect 433352 26206 434116 26234
rect 431960 24608 432012 24614
rect 431960 24550 432012 24556
rect 430580 21888 430632 21894
rect 430580 21830 430632 21836
rect 430580 21616 430632 21622
rect 430580 21558 430632 21564
rect 430592 16574 430620 21558
rect 432064 17746 432092 26206
rect 432144 24744 432196 24750
rect 432144 24686 432196 24692
rect 432052 17740 432104 17746
rect 432052 17682 432104 17688
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 432156 6914 432184 24686
rect 433352 15094 433380 26206
rect 434824 23322 434852 29786
rect 435008 26994 435036 29838
rect 435927 29786 435979 29792
rect 436204 29838 436885 29866
rect 437768 29838 437803 29866
rect 438596 29838 438704 29866
rect 439516 29838 439622 29866
rect 440436 29838 440523 29866
rect 440712 29838 441441 29866
rect 441632 29838 442359 29866
rect 443012 29838 443209 29866
rect 443288 29838 444161 29866
rect 444944 29838 445062 29866
rect 445772 29838 445963 29866
rect 446232 29838 446881 29866
rect 447152 29838 447782 29866
rect 448520 29844 448572 29850
rect 434996 26988 435048 26994
rect 434996 26930 435048 26936
rect 436100 26988 436152 26994
rect 436100 26930 436152 26936
rect 434812 23316 434864 23322
rect 434812 23258 434864 23264
rect 434720 20460 434772 20466
rect 434720 20402 434772 20408
rect 434732 16574 434760 20402
rect 434732 16546 435128 16574
rect 433340 15088 433392 15094
rect 433340 15030 433392 15036
rect 434444 8356 434496 8362
rect 434444 8298 434496 8304
rect 432064 6886 432184 6914
rect 432064 480 432092 6886
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 434456 480 434484 8298
rect 429630 354 429742 480
rect 429396 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 436112 6914 436140 26930
rect 436204 16522 436232 29838
rect 437768 27130 437796 29838
rect 437756 27124 437808 27130
rect 437756 27066 437808 27072
rect 438596 26234 438624 29838
rect 439516 26234 439544 29838
rect 440436 27198 440464 29838
rect 440424 27192 440476 27198
rect 440424 27134 440476 27140
rect 440240 27056 440292 27062
rect 440240 26998 440292 27004
rect 437584 26206 438624 26234
rect 438872 26206 439544 26234
rect 437584 19038 437612 26206
rect 437572 19032 437624 19038
rect 437572 18974 437624 18980
rect 436192 16516 436244 16522
rect 436192 16458 436244 16464
rect 438872 13054 438900 26206
rect 439136 13728 439188 13734
rect 439136 13670 439188 13676
rect 438860 13048 438912 13054
rect 438860 12990 438912 12996
rect 437940 8968 437992 8974
rect 437940 8910 437992 8916
rect 436112 6886 436784 6914
rect 436756 480 436784 6886
rect 437952 480 437980 8910
rect 439148 480 439176 13670
rect 440252 3074 440280 26998
rect 440712 26234 440740 29838
rect 440436 26206 440740 26234
rect 440332 25764 440384 25770
rect 440332 25706 440384 25712
rect 440344 3262 440372 25706
rect 440436 22030 440464 26206
rect 441632 26110 441660 29838
rect 441620 26104 441672 26110
rect 441620 26046 441672 26052
rect 440424 22024 440476 22030
rect 440424 21966 440476 21972
rect 441620 19168 441672 19174
rect 441620 19110 441672 19116
rect 441632 16574 441660 19110
rect 441632 16546 442672 16574
rect 440332 3256 440384 3262
rect 440332 3198 440384 3204
rect 441528 3256 441580 3262
rect 441528 3198 441580 3204
rect 440252 3046 440372 3074
rect 440344 480 440372 3046
rect 441540 480 441568 3198
rect 442644 480 442672 16546
rect 443012 10878 443040 29838
rect 443288 26234 443316 29838
rect 444944 26234 444972 29838
rect 443104 26206 443316 26234
rect 444392 26206 444972 26234
rect 443104 15162 443132 26206
rect 443092 15156 443144 15162
rect 443092 15098 443144 15104
rect 443000 10872 443052 10878
rect 443000 10814 443052 10820
rect 444392 9586 444420 26206
rect 445772 10810 445800 29838
rect 446232 26234 446260 29838
rect 445864 26206 446260 26234
rect 445864 14618 445892 26206
rect 447152 24410 447180 29838
rect 448520 29786 448572 29792
rect 448624 29838 448717 29866
rect 449590 29850 449618 30049
rect 450508 29866 450536 30049
rect 451409 29866 451437 30049
rect 452327 29866 452355 30049
rect 453228 29866 453256 30049
rect 454163 29866 454191 30049
rect 455013 29866 455041 30049
rect 455965 29866 455993 30049
rect 449578 29844 449630 29850
rect 447232 27124 447284 27130
rect 447232 27066 447284 27072
rect 447140 24404 447192 24410
rect 447140 24346 447192 24352
rect 447244 16574 447272 27066
rect 447244 16546 447456 16574
rect 445852 14612 445904 14618
rect 445852 14554 445904 14560
rect 445852 12300 445904 12306
rect 445852 12242 445904 12248
rect 445760 10804 445812 10810
rect 445760 10746 445812 10752
rect 444380 9580 444432 9586
rect 444380 9522 444432 9528
rect 445024 5160 445076 5166
rect 445024 5102 445076 5108
rect 443828 3256 443880 3262
rect 443828 3198 443880 3204
rect 443840 480 443868 3198
rect 445036 480 445064 5102
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445864 354 445892 12242
rect 447428 480 447456 16546
rect 448532 3369 448560 29786
rect 448624 16590 448652 29838
rect 449578 29786 449630 29792
rect 450464 29838 450536 29866
rect 451292 29838 451437 29866
rect 452304 29838 452355 29866
rect 453224 29838 453256 29866
rect 454144 29838 454191 29866
rect 454236 29838 455041 29866
rect 455432 29838 455993 29866
rect 456849 29866 456877 30049
rect 457767 29866 457795 30049
rect 458668 29866 458696 30049
rect 456849 29838 456932 29866
rect 449900 27192 449952 27198
rect 449900 27134 449952 27140
rect 448796 17468 448848 17474
rect 448796 17410 448848 17416
rect 448612 16584 448664 16590
rect 448612 16526 448664 16532
rect 448704 12232 448756 12238
rect 448704 12174 448756 12180
rect 448612 4208 448664 4214
rect 448612 4150 448664 4156
rect 448624 3738 448652 4150
rect 448716 3738 448744 12174
rect 448612 3732 448664 3738
rect 448612 3674 448664 3680
rect 448704 3732 448756 3738
rect 448704 3674 448756 3680
rect 448808 3482 448836 17410
rect 449808 3732 449860 3738
rect 449808 3674 449860 3680
rect 448624 3454 448836 3482
rect 448518 3360 448574 3369
rect 448518 3295 448574 3304
rect 448624 480 448652 3454
rect 449820 480 449848 3674
rect 449912 3482 449940 27134
rect 450464 26234 450492 29838
rect 450004 26206 450492 26234
rect 450004 4214 450032 26206
rect 449992 4208 450044 4214
rect 449992 4150 450044 4156
rect 449912 3454 450952 3482
rect 451292 3466 451320 29838
rect 452304 26234 452332 29838
rect 453224 26234 453252 29838
rect 454040 27328 454092 27334
rect 454040 27270 454092 27276
rect 453304 27260 453356 27266
rect 453304 27202 453356 27208
rect 451384 26206 452332 26234
rect 452672 26206 453252 26234
rect 451384 3534 451412 26206
rect 451648 13320 451700 13326
rect 451648 13262 451700 13268
rect 451372 3528 451424 3534
rect 451372 3470 451424 3476
rect 450924 480 450952 3454
rect 451280 3460 451332 3466
rect 451280 3402 451332 3408
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 13262
rect 452672 3602 452700 26206
rect 453316 16574 453344 27202
rect 453316 16546 453436 16574
rect 453304 12164 453356 12170
rect 453304 12106 453356 12112
rect 452660 3596 452712 3602
rect 452660 3538 452712 3544
rect 453316 480 453344 12106
rect 453408 11762 453436 16546
rect 453396 11756 453448 11762
rect 453396 11698 453448 11704
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 27270
rect 454144 3670 454172 29838
rect 454236 3806 454264 29838
rect 455432 3874 455460 29838
rect 456800 28144 456852 28150
rect 456800 28086 456852 28092
rect 455512 20188 455564 20194
rect 455512 20130 455564 20136
rect 455524 16574 455552 20130
rect 455524 16546 455736 16574
rect 455420 3868 455472 3874
rect 455420 3810 455472 3816
rect 454224 3800 454276 3806
rect 454224 3742 454276 3748
rect 454132 3664 454184 3670
rect 454132 3606 454184 3612
rect 455708 480 455736 16546
rect 456812 4010 456840 28086
rect 456904 16574 456932 29838
rect 457732 29838 457795 29866
rect 458652 29838 458696 29866
rect 459586 29866 459614 30049
rect 460504 29866 460532 30049
rect 461422 29866 461450 30049
rect 459586 29838 459692 29866
rect 457732 28150 457760 29838
rect 457720 28144 457772 28150
rect 457720 28086 457772 28092
rect 458652 26234 458680 29838
rect 459560 28144 459612 28150
rect 459560 28086 459612 28092
rect 458192 26206 458680 26234
rect 456904 16546 457024 16574
rect 456800 4004 456852 4010
rect 456800 3946 456852 3952
rect 456996 3942 457024 16546
rect 457076 12096 457128 12102
rect 457076 12038 457128 12044
rect 456984 3936 457036 3942
rect 456984 3878 457036 3884
rect 457088 3482 457116 12038
rect 458192 4078 458220 26206
rect 458272 24268 458324 24274
rect 458272 24210 458324 24216
rect 458284 16574 458312 24210
rect 458284 16546 459232 16574
rect 458180 4072 458232 4078
rect 458180 4014 458232 4020
rect 456904 3454 457116 3482
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 456904 480 456932 3454
rect 458100 480 458128 3470
rect 459204 480 459232 16546
rect 459572 3398 459600 28086
rect 459664 4146 459692 29838
rect 460492 29838 460532 29866
rect 461412 29838 461450 29866
rect 462323 29866 462351 30049
rect 463241 29866 463269 30049
rect 464159 29866 464187 30049
rect 465060 29866 465088 30049
rect 465978 29866 466006 30049
rect 466828 29866 466856 30049
rect 467763 29866 467791 30049
rect 468681 29866 468709 30049
rect 462323 29838 462360 29866
rect 463241 29838 463280 29866
rect 464159 29838 464200 29866
rect 465060 29838 465120 29866
rect 465978 29838 466040 29866
rect 466828 29838 466868 29866
rect 460492 28150 460520 29838
rect 460480 28144 460532 28150
rect 460480 28086 460532 28092
rect 461032 27532 461084 27538
rect 461032 27474 461084 27480
rect 461044 16574 461072 27474
rect 461412 26926 461440 29838
rect 461400 26920 461452 26926
rect 461400 26862 461452 26868
rect 462332 26234 462360 29838
rect 463252 26994 463280 29838
rect 464172 27062 464200 29838
rect 464160 27056 464212 27062
rect 464160 26998 464212 27004
rect 463240 26988 463292 26994
rect 463240 26930 463292 26936
rect 465092 26234 465120 29838
rect 465264 27600 465316 27606
rect 465264 27542 465316 27548
rect 462332 26206 462544 26234
rect 465092 26206 465212 26234
rect 462412 18828 462464 18834
rect 462412 18770 462464 18776
rect 461044 16546 461624 16574
rect 459928 12028 459980 12034
rect 459928 11970 459980 11976
rect 459652 4140 459704 4146
rect 459652 4082 459704 4088
rect 459560 3392 459612 3398
rect 459560 3334 459612 3340
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 11970
rect 461596 480 461624 16546
rect 461676 16448 461728 16454
rect 461676 16390 461728 16396
rect 461688 3466 461716 16390
rect 461676 3460 461728 3466
rect 461676 3402 461728 3408
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 18770
rect 462516 3330 462544 26206
rect 464344 25900 464396 25906
rect 464344 25842 464396 25848
rect 463976 11960 464028 11966
rect 463976 11902 464028 11908
rect 462504 3324 462556 3330
rect 462504 3266 462556 3272
rect 463988 480 464016 11902
rect 464356 3602 464384 25842
rect 465184 16574 465212 26206
rect 465092 16546 465212 16574
rect 464344 3596 464396 3602
rect 464344 3538 464396 3544
rect 465092 3262 465120 16546
rect 465276 6914 465304 27542
rect 466012 27130 466040 29838
rect 466840 27198 466868 29838
rect 467760 29838 467791 29866
rect 467944 29838 468709 29866
rect 469582 29866 469610 30049
rect 470500 29866 470528 30049
rect 471401 29866 471429 30049
rect 472336 29866 472364 30049
rect 469582 29838 469628 29866
rect 470500 29838 470548 29866
rect 467760 27334 467788 29838
rect 467748 27328 467800 27334
rect 467748 27270 467800 27276
rect 466828 27192 466880 27198
rect 466828 27134 466880 27140
rect 466000 27124 466052 27130
rect 466000 27066 466052 27072
rect 467840 26308 467892 26314
rect 467840 26250 467892 26256
rect 466460 23248 466512 23254
rect 466460 23190 466512 23196
rect 466472 16574 466500 23190
rect 466472 16546 467512 16574
rect 465184 6886 465304 6914
rect 465080 3256 465132 3262
rect 465080 3198 465132 3204
rect 465184 480 465212 6886
rect 466276 2100 466328 2106
rect 466276 2042 466328 2048
rect 466288 480 466316 2042
rect 467484 480 467512 16546
rect 467852 490 467880 26250
rect 467944 3534 467972 29838
rect 469600 27538 469628 29838
rect 470520 27606 470548 29838
rect 471348 29838 471429 29866
rect 472268 29838 472364 29866
rect 473237 29866 473265 30049
rect 474155 29866 474183 30049
rect 475056 29866 475084 30049
rect 473237 29838 473308 29866
rect 470508 27600 470560 27606
rect 470508 27542 470560 27548
rect 469588 27532 469640 27538
rect 469588 27474 469640 27480
rect 471348 26314 471376 29838
rect 471336 26308 471388 26314
rect 471336 26250 471388 26256
rect 472268 26234 472296 29838
rect 473280 27606 473308 29838
rect 473372 29838 474183 29866
rect 474832 29844 474884 29850
rect 473268 27600 473320 27606
rect 473268 27542 473320 27548
rect 471992 26206 472296 26234
rect 471992 16574 472020 26206
rect 471992 16546 472296 16574
rect 469864 10396 469916 10402
rect 469864 10338 469916 10344
rect 467932 3528 467984 3534
rect 467932 3470 467984 3476
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 467852 462 468248 490
rect 469876 480 469904 10338
rect 471060 9512 471112 9518
rect 471060 9454 471112 9460
rect 471072 480 471100 9454
rect 472268 480 472296 16546
rect 473372 3058 473400 29838
rect 474832 29786 474884 29792
rect 475028 29838 475084 29866
rect 475991 29850 476019 30049
rect 476875 29866 476903 30049
rect 477810 29866 477838 30049
rect 475979 29844 476031 29850
rect 474740 27600 474792 27606
rect 474740 27542 474792 27548
rect 473452 15972 473504 15978
rect 473452 15914 473504 15920
rect 473360 3052 473412 3058
rect 473360 2994 473412 3000
rect 473464 480 473492 15914
rect 474556 3596 474608 3602
rect 474556 3538 474608 3544
rect 474568 480 474596 3538
rect 474752 3482 474780 27542
rect 474844 3602 474872 29786
rect 475028 26234 475056 29838
rect 475979 29786 476031 29792
rect 476132 29838 476903 29866
rect 477788 29838 477838 29866
rect 478660 29866 478688 30049
rect 479595 29866 479623 30049
rect 480496 29866 480524 30049
rect 481414 29866 481442 30049
rect 482315 29866 482343 30049
rect 483250 29866 483278 30049
rect 484151 29866 484179 30049
rect 485069 29866 485097 30049
rect 478660 29838 478736 29866
rect 474936 26206 475056 26234
rect 474936 3670 474964 26206
rect 474924 3664 474976 3670
rect 474924 3606 474976 3612
rect 474832 3596 474884 3602
rect 474832 3538 474884 3544
rect 476132 3534 476160 29838
rect 477788 26926 477816 29838
rect 477776 26920 477828 26926
rect 477776 26862 477828 26868
rect 478708 26314 478736 29838
rect 478892 29838 479623 29866
rect 480456 29838 480524 29866
rect 481376 29838 481442 29866
rect 482296 29838 482343 29866
rect 483032 29838 483278 29866
rect 483584 29838 484179 29866
rect 484412 29838 485097 29866
rect 485970 29866 485998 30049
rect 486888 29866 486916 30049
rect 487806 29866 487834 30049
rect 488690 29866 488718 30049
rect 485970 29838 486004 29866
rect 478696 26308 478748 26314
rect 478696 26250 478748 26256
rect 478892 10402 478920 29838
rect 480456 27130 480484 29838
rect 481376 27606 481404 29838
rect 481364 27600 481416 27606
rect 481364 27542 481416 27548
rect 480444 27124 480496 27130
rect 480444 27066 480496 27072
rect 482296 26994 482324 29838
rect 482284 26988 482336 26994
rect 482284 26930 482336 26936
rect 482284 26308 482336 26314
rect 482284 26250 482336 26256
rect 478880 10396 478932 10402
rect 478880 10338 478932 10344
rect 476488 10328 476540 10334
rect 476488 10270 476540 10276
rect 476120 3528 476172 3534
rect 474752 3454 475792 3482
rect 476120 3470 476172 3476
rect 475764 480 475792 3454
rect 468220 354 468248 462
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 10270
rect 482296 9042 482324 26250
rect 480536 9036 480588 9042
rect 480536 8978 480588 8984
rect 482284 9036 482336 9042
rect 482284 8978 482336 8984
rect 478144 3460 478196 3466
rect 478144 3402 478196 3408
rect 478156 480 478184 3402
rect 479340 3052 479392 3058
rect 479340 2994 479392 3000
rect 479352 480 479380 2994
rect 480548 480 480576 8978
rect 483032 8974 483060 29838
rect 483584 26234 483612 29838
rect 483124 26206 483612 26234
rect 483124 10334 483152 26206
rect 483204 17400 483256 17406
rect 483204 17342 483256 17348
rect 483216 16574 483244 17342
rect 483216 16546 484072 16574
rect 483112 10328 483164 10334
rect 483112 10270 483164 10276
rect 483020 8968 483072 8974
rect 483020 8910 483072 8916
rect 481732 6656 481784 6662
rect 481732 6598 481784 6604
rect 481744 480 481772 6598
rect 482836 3664 482888 3670
rect 482836 3606 482888 3612
rect 482848 480 482876 3606
rect 484044 480 484072 16546
rect 484412 11830 484440 29838
rect 485044 27600 485096 27606
rect 485044 27542 485096 27548
rect 485056 11898 485084 27542
rect 485976 27062 486004 29838
rect 486804 29838 486916 29866
rect 487724 29838 487834 29866
rect 488540 29844 488592 29850
rect 485964 27056 486016 27062
rect 485964 26998 486016 27004
rect 486804 26234 486832 29838
rect 487724 26234 487752 29838
rect 488540 29786 488592 29792
rect 488644 29838 488718 29866
rect 489625 29850 489653 30049
rect 489613 29844 489665 29850
rect 485792 26206 486832 26234
rect 487264 26206 487752 26234
rect 485792 13190 485820 26206
rect 487264 18766 487292 26206
rect 487160 18760 487212 18766
rect 487160 18702 487212 18708
rect 487252 18760 487304 18766
rect 487252 18702 487304 18708
rect 485780 13184 485832 13190
rect 485780 13126 485832 13132
rect 485044 11892 485096 11898
rect 485044 11834 485096 11840
rect 484400 11824 484452 11830
rect 484400 11766 484452 11772
rect 485228 6588 485280 6594
rect 485228 6530 485280 6536
rect 485240 480 485268 6530
rect 486424 3596 486476 3602
rect 486424 3538 486476 3544
rect 486436 480 486464 3538
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 18702
rect 488552 3262 488580 29786
rect 488644 15978 488672 29838
rect 490526 29832 490554 30049
rect 489613 29786 489665 29792
rect 490484 29804 490554 29832
rect 491300 29844 491352 29850
rect 490484 26234 490512 29804
rect 491410 29832 491438 30049
rect 492328 29850 492356 30049
rect 491300 29786 491352 29792
rect 491404 29804 491438 29832
rect 492316 29844 492368 29850
rect 489932 26206 490512 26234
rect 488632 15972 488684 15978
rect 488632 15914 488684 15920
rect 489932 6914 489960 26206
rect 490012 21548 490064 21554
rect 490012 21490 490064 21496
rect 490024 16574 490052 21490
rect 490024 16546 490696 16574
rect 489932 6886 490052 6914
rect 488816 6520 488868 6526
rect 488816 6462 488868 6468
rect 488540 3256 488592 3262
rect 488540 3198 488592 3204
rect 488828 480 488856 6462
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 489932 480 489960 3470
rect 490024 3330 490052 6886
rect 490012 3324 490064 3330
rect 490012 3266 490064 3272
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 491312 4146 491340 29786
rect 491300 4140 491352 4146
rect 491300 4082 491352 4088
rect 491404 3398 491432 29804
rect 493229 29832 493257 30049
rect 492316 29786 492368 29792
rect 492784 29804 493257 29832
rect 494060 29844 494112 29850
rect 492680 26920 492732 26926
rect 492680 26862 492732 26868
rect 492312 13592 492364 13598
rect 492312 13534 492364 13540
rect 491392 3392 491444 3398
rect 491392 3334 491444 3340
rect 492324 480 492352 13534
rect 492692 490 492720 26862
rect 492784 4078 492812 29804
rect 494147 29832 494175 30049
rect 495065 29850 495093 30049
rect 495053 29844 495105 29850
rect 494147 29804 494192 29832
rect 494060 29786 494112 29792
rect 492772 4072 492824 4078
rect 492772 4014 492824 4020
rect 494072 3942 494100 29786
rect 494164 4010 494192 29804
rect 495983 29832 496011 30049
rect 496884 29832 496912 30049
rect 497802 29832 497830 30049
rect 498703 29832 498731 30049
rect 499638 29866 499666 30049
rect 500505 29866 500533 30049
rect 501457 29866 501485 30049
rect 499638 29838 499712 29866
rect 500505 29838 500540 29866
rect 495053 29786 495105 29792
rect 495452 29804 496011 29832
rect 496832 29804 496912 29832
rect 497752 29804 497830 29832
rect 498396 29804 498731 29832
rect 494244 20120 494296 20126
rect 494244 20062 494296 20068
rect 494256 16574 494284 20062
rect 494256 16546 494744 16574
rect 494152 4004 494204 4010
rect 494152 3946 494204 3952
rect 494060 3936 494112 3942
rect 494060 3878 494112 3884
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 492692 462 493088 490
rect 494716 480 494744 16546
rect 495452 3874 495480 29804
rect 495532 14544 495584 14550
rect 495532 14486 495584 14492
rect 495440 3868 495492 3874
rect 495440 3810 495492 3816
rect 493060 354 493088 462
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495544 354 495572 14486
rect 496832 3806 496860 29804
rect 497752 26234 497780 29804
rect 496924 26206 497780 26234
rect 496820 3800 496872 3806
rect 496820 3742 496872 3748
rect 496924 3738 496952 26206
rect 498292 22908 498344 22914
rect 498292 22850 498344 22856
rect 497096 9036 497148 9042
rect 497096 8978 497148 8984
rect 496912 3732 496964 3738
rect 496912 3674 496964 3680
rect 497108 480 497136 8978
rect 498304 6914 498332 22850
rect 498212 6886 498332 6914
rect 498212 480 498240 6886
rect 498396 3670 498424 29804
rect 499580 10396 499632 10402
rect 499580 10338 499632 10344
rect 499396 6452 499448 6458
rect 499396 6394 499448 6400
rect 498384 3664 498436 3670
rect 498384 3606 498436 3612
rect 499408 480 499436 6394
rect 499592 3482 499620 10338
rect 499684 3602 499712 29838
rect 500512 26926 500540 29838
rect 500972 29838 501485 29866
rect 502324 29866 502352 30049
rect 502885 29866 502913 30048
rect 502324 29838 502380 29866
rect 500500 26920 500552 26926
rect 500500 26862 500552 26868
rect 499672 3596 499724 3602
rect 499672 3538 499724 3544
rect 499592 3454 500632 3482
rect 500972 3466 501000 29838
rect 501052 25696 501104 25702
rect 501052 25638 501104 25644
rect 501064 16574 501092 25638
rect 501064 16546 501368 16574
rect 500604 480 500632 3454
rect 500960 3460 501012 3466
rect 500960 3402 501012 3408
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502352 3602 502380 29838
rect 502444 29838 502913 29866
rect 502340 3596 502392 3602
rect 502340 3538 502392 3544
rect 502444 3369 502472 29838
rect 503720 27124 503772 27130
rect 503720 27066 503772 27072
rect 502984 6384 503036 6390
rect 502984 6326 503036 6332
rect 502430 3360 502486 3369
rect 502430 3295 502486 3304
rect 502996 480 503024 6326
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 27066
rect 512644 27056 512696 27062
rect 512644 26998 512696 27004
rect 510620 26988 510672 26994
rect 510620 26930 510672 26936
rect 505100 24200 505152 24206
rect 505100 24142 505152 24148
rect 505112 16574 505140 24142
rect 510632 16574 510660 26930
rect 505112 16546 505416 16574
rect 510632 16546 511304 16574
rect 505388 480 505416 16546
rect 508872 13116 508924 13122
rect 508872 13058 508924 13064
rect 507216 11892 507268 11898
rect 507216 11834 507268 11840
rect 506480 6316 506532 6322
rect 506480 6258 506532 6264
rect 506492 480 506520 6258
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 11834
rect 508884 480 508912 13058
rect 510068 6248 510120 6254
rect 510068 6190 510120 6196
rect 510080 480 510108 6190
rect 511276 480 511304 16546
rect 512656 6254 512684 26998
rect 569224 26920 569276 26926
rect 569224 26862 569276 26868
rect 547880 25628 547932 25634
rect 547880 25570 547932 25576
rect 516140 24472 516192 24478
rect 516140 24414 516192 24420
rect 514760 17332 514812 17338
rect 514760 17274 514812 17280
rect 514772 16574 514800 17274
rect 516152 16574 516180 24414
rect 534080 23044 534132 23050
rect 534080 22986 534132 22992
rect 529940 22840 529992 22846
rect 529940 22782 529992 22788
rect 523040 21480 523092 21486
rect 523040 21422 523092 21428
rect 518900 18692 518952 18698
rect 518900 18634 518952 18640
rect 518912 16574 518940 18634
rect 514772 16546 515536 16574
rect 516152 16546 517192 16574
rect 518912 16546 519584 16574
rect 514760 8968 514812 8974
rect 514760 8910 514812 8916
rect 512644 6248 512696 6254
rect 512644 6190 512696 6196
rect 513564 6180 513616 6186
rect 513564 6122 513616 6128
rect 512460 5092 512512 5098
rect 512460 5034 512512 5040
rect 512472 480 512500 5034
rect 513576 480 513604 6122
rect 514772 480 514800 8910
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517164 480 517192 16546
rect 517888 10328 517940 10334
rect 517888 10270 517940 10276
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 10270
rect 519556 480 519584 16546
rect 520280 15904 520332 15910
rect 520280 15846 520332 15852
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 15846
rect 521660 11824 521712 11830
rect 521660 11766 521712 11772
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 11766
rect 523052 480 523080 21422
rect 525800 20052 525852 20058
rect 525800 19994 525852 20000
rect 525812 16574 525840 19994
rect 525812 16546 526208 16574
rect 524236 9376 524288 9382
rect 524236 9318 524288 9324
rect 524248 480 524276 9318
rect 525432 6248 525484 6254
rect 525432 6190 525484 6196
rect 525444 480 525472 6190
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 13456 527876 13462
rect 527824 13398 527876 13404
rect 527836 480 527864 13398
rect 528560 13184 528612 13190
rect 528560 13126 528612 13132
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 13126
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 22782
rect 531320 18760 531372 18766
rect 531320 18702 531372 18708
rect 531332 3194 531360 18702
rect 534092 16574 534120 22986
rect 538220 21684 538272 21690
rect 538220 21626 538272 21632
rect 534092 16546 534488 16574
rect 531412 10464 531464 10470
rect 531412 10406 531464 10412
rect 531320 3188 531372 3194
rect 531320 3130 531372 3136
rect 531424 3074 531452 10406
rect 533712 5024 533764 5030
rect 533712 4966 533764 4972
rect 532148 3188 532200 3194
rect 532148 3130 532200 3136
rect 531332 3046 531452 3074
rect 531332 480 531360 3046
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3130
rect 533724 480 533752 4966
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536104 15972 536156 15978
rect 536104 15914 536156 15920
rect 536116 480 536144 15914
rect 537208 4956 537260 4962
rect 537208 4898 537260 4904
rect 537220 480 537248 4898
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 21626
rect 540980 17672 541032 17678
rect 540980 17614 541032 17620
rect 540992 16574 541020 17614
rect 540992 16546 542032 16574
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 539600 3256 539652 3262
rect 539600 3198 539652 3204
rect 539612 480 539640 3198
rect 540808 480 540836 4830
rect 542004 480 542032 16546
rect 545488 16108 545540 16114
rect 545488 16050 545540 16056
rect 544384 4820 544436 4826
rect 544384 4762 544436 4768
rect 543188 3324 543240 3330
rect 543188 3266 543240 3272
rect 543200 480 543228 3266
rect 544396 480 544424 4762
rect 545500 480 545528 16050
rect 546684 3392 546736 3398
rect 546684 3334 546736 3340
rect 546696 480 546724 3334
rect 547892 480 547920 25570
rect 550640 24132 550692 24138
rect 550640 24074 550692 24080
rect 550652 16574 550680 24074
rect 564532 21412 564584 21418
rect 564532 21354 564584 21360
rect 561680 18624 561732 18630
rect 561680 18566 561732 18572
rect 557540 17264 557592 17270
rect 557540 17206 557592 17212
rect 557552 16574 557580 17206
rect 561692 16574 561720 18566
rect 564544 16574 564572 21354
rect 568580 19984 568632 19990
rect 568580 19926 568632 19932
rect 568592 16574 568620 19926
rect 550652 16546 551048 16574
rect 557552 16546 558592 16574
rect 561692 16546 562088 16574
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 549076 8084 549128 8090
rect 549076 8026 549128 8032
rect 549088 480 549116 8026
rect 550272 4140 550324 4146
rect 550272 4082 550324 4088
rect 550284 480 550312 4082
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 554780 14476 554832 14482
rect 554780 14418 554832 14424
rect 552664 8016 552716 8022
rect 552664 7958 552716 7964
rect 552676 480 552704 7958
rect 553768 4072 553820 4078
rect 553768 4014 553820 4020
rect 553780 480 553808 4014
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 14418
rect 556160 7948 556212 7954
rect 556160 7890 556212 7896
rect 556172 480 556200 7890
rect 557356 4004 557408 4010
rect 557356 3946 557408 3952
rect 557368 480 557396 3946
rect 558564 480 558592 16546
rect 559748 7880 559800 7886
rect 559748 7822 559800 7828
rect 559760 480 559788 7822
rect 560852 3936 560904 3942
rect 560852 3878 560904 3884
rect 560864 480 560892 3878
rect 562060 480 562088 16546
rect 563060 14884 563112 14890
rect 563060 14826 563112 14832
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 14826
rect 564440 3868 564492 3874
rect 564440 3810 564492 3816
rect 564452 480 564480 3810
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566832 11756 566884 11762
rect 566832 11698 566884 11704
rect 566844 480 566872 11698
rect 568028 3800 568080 3806
rect 568028 3742 568080 3748
rect 568040 480 568068 3742
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 16546
rect 569236 4826 569264 26862
rect 575480 25560 575532 25566
rect 575480 25502 575532 25508
rect 572720 22772 572772 22778
rect 572720 22714 572772 22720
rect 570328 7812 570380 7818
rect 570328 7754 570380 7760
rect 569224 4820 569276 4826
rect 569224 4762 569276 4768
rect 570340 480 570368 7754
rect 571524 3732 571576 3738
rect 571524 3674 571576 3680
rect 571536 480 571564 3674
rect 572732 480 572760 22714
rect 575492 16574 575520 25502
rect 575492 16546 575888 16574
rect 573916 7744 573968 7750
rect 573916 7686 573968 7692
rect 573928 480 573956 7686
rect 575112 3664 575164 3670
rect 575112 3606 575164 3612
rect 575124 480 575152 3606
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 7676 577464 7682
rect 577412 7618 577464 7624
rect 577424 480 577452 7618
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 578620 480 578648 3470
rect 579816 480 579844 4762
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 6458 3304 6514 3360
rect 150530 3576 150586 3632
rect 383566 3304 383622 3360
rect 448518 3304 448574 3360
rect 502430 3304 502486 3360
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 150525 3634 150591 3637
rect 137970 3632 150591 3634
rect 137970 3576 150530 3632
rect 150586 3576 150591 3632
rect 137970 3574 150591 3576
rect 6453 3362 6519 3365
rect 137970 3362 138030 3574
rect 150525 3571 150591 3574
rect 6453 3360 138030 3362
rect 6453 3304 6458 3360
rect 6514 3304 138030 3360
rect 6453 3302 138030 3304
rect 383561 3362 383627 3365
rect 448513 3362 448579 3365
rect 383561 3360 448579 3362
rect 383561 3304 383566 3360
rect 383622 3304 448518 3360
rect 448574 3304 448579 3360
rect 383561 3302 448579 3304
rect 6453 3299 6519 3302
rect 383561 3299 383627 3302
rect 448513 3299 448579 3302
rect 502425 3362 502491 3365
rect 583385 3362 583451 3365
rect 502425 3360 583451 3362
rect 502425 3304 502430 3360
rect 502486 3304 583390 3360
rect 583446 3304 583451 3360
rect 502425 3302 583451 3304
rect 502425 3299 502491 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 475836 56414 488898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 475836 60134 492618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 475836 63854 496338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 475836 67574 500058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 475836 74414 506898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475836 78134 510618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 475836 81854 478338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 475836 85574 482058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 475836 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 475836 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 475836 99854 496338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 475836 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 475836 110414 506898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475836 114134 510618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 475836 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 475836 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 475836 128414 488898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 475836 132134 492618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 475836 135854 496338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 475836 139574 500058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 475836 146414 506898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475836 150134 510618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 475836 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 475836 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 475836 164414 488898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 475836 168134 492618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 475836 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 475836 175574 500058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 475836 182414 506898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475836 186134 510618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 475836 189854 478338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 475836 193574 482058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 475836 200414 488898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 475836 204134 492618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 475836 207854 496338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 475836 211574 500058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 475836 218414 506898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475836 222134 510618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 475836 225854 478338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 475836 229574 482058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 475836 236414 488898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 475836 240134 492618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 475836 243854 496338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 475836 247574 500058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 475836 254414 506898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475836 258134 510618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 475836 261854 478338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 475836 265574 482058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 475836 272414 488898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 475836 276134 492618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 475836 279854 496338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 475836 283574 500058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 475836 290414 506898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475836 294134 510618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 475836 297854 478338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 475836 301574 482058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 475836 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 475836 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 475836 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 475836 319574 500058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 475836 326414 506898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475836 330134 510618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 475836 333854 478338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 475836 337574 482058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 475836 344414 488898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 475836 348134 492618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 475836 351854 496338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 475836 355574 500058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 475836 362414 506898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475836 366134 510618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 475836 369854 478338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 475836 373574 482058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 475836 380414 488898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 475836 384134 492618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 475836 387854 496338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 475836 391574 500058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 475836 398414 506898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475836 402134 510618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 475836 405854 478338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 475836 409574 482058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 475836 416414 488898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 475836 420134 492618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 475836 423854 496338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 475836 427574 500058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 475836 434414 506898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475836 438134 510618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 475836 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 475836 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 475836 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 475836 456134 492618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 475836 459854 496338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 475836 463574 500058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 475836 470414 506898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475836 474134 510618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 475836 477854 478338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 475836 481574 482058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 475836 488414 488898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 475836 492134 492618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 475836 495854 496338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 475836 499574 500058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 475836 506414 506898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475836 510134 510618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 475836 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 475836 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 58960 453454 61960 453486
rect 58960 453218 59062 453454
rect 59298 453218 59382 453454
rect 59618 453218 59702 453454
rect 59938 453218 60022 453454
rect 60258 453218 60342 453454
rect 60578 453218 60662 453454
rect 60898 453218 60982 453454
rect 61218 453218 61302 453454
rect 61538 453218 61622 453454
rect 61858 453218 61960 453454
rect 58960 453134 61960 453218
rect 58960 452898 59062 453134
rect 59298 452898 59382 453134
rect 59618 452898 59702 453134
rect 59938 452898 60022 453134
rect 60258 452898 60342 453134
rect 60578 452898 60662 453134
rect 60898 452898 60982 453134
rect 61218 452898 61302 453134
rect 61538 452898 61622 453134
rect 61858 452898 61960 453134
rect 58960 452866 61960 452898
rect 71121 453454 71469 453486
rect 71121 453218 71177 453454
rect 71413 453218 71469 453454
rect 71121 453134 71469 453218
rect 71121 452898 71177 453134
rect 71413 452898 71469 453134
rect 71121 452866 71469 452898
rect 166185 453454 166533 453486
rect 166185 453218 166241 453454
rect 166477 453218 166533 453454
rect 166185 453134 166533 453218
rect 166185 452898 166241 453134
rect 166477 452898 166533 453134
rect 166185 452866 166533 452898
rect 403077 453454 403425 453486
rect 403077 453218 403133 453454
rect 403369 453218 403425 453454
rect 403077 453134 403425 453218
rect 403077 452898 403133 453134
rect 403369 452898 403425 453134
rect 403077 452866 403425 452898
rect 498141 453454 498489 453486
rect 498141 453218 498197 453454
rect 498433 453218 498489 453454
rect 498141 453134 498489 453218
rect 498141 452898 498197 453134
rect 498433 452898 498489 453134
rect 498141 452866 498489 452898
rect 507948 453454 510948 453486
rect 507948 453218 508050 453454
rect 508286 453218 508370 453454
rect 508606 453218 508690 453454
rect 508926 453218 509010 453454
rect 509246 453218 509330 453454
rect 509566 453218 509650 453454
rect 509886 453218 509970 453454
rect 510206 453218 510290 453454
rect 510526 453218 510610 453454
rect 510846 453218 510948 453454
rect 507948 453134 510948 453218
rect 507948 452898 508050 453134
rect 508286 452898 508370 453134
rect 508606 452898 508690 453134
rect 508926 452898 509010 453134
rect 509246 452898 509330 453134
rect 509566 452898 509650 453134
rect 509886 452898 509970 453134
rect 510206 452898 510290 453134
rect 510526 452898 510610 453134
rect 510846 452898 510948 453134
rect 507948 452866 510948 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 62960 435454 65960 435486
rect 62960 435218 63062 435454
rect 63298 435218 63382 435454
rect 63618 435218 63702 435454
rect 63938 435218 64022 435454
rect 64258 435218 64342 435454
rect 64578 435218 64662 435454
rect 64898 435218 64982 435454
rect 65218 435218 65302 435454
rect 65538 435218 65622 435454
rect 65858 435218 65960 435454
rect 62960 435134 65960 435218
rect 62960 434898 63062 435134
rect 63298 434898 63382 435134
rect 63618 434898 63702 435134
rect 63938 434898 64022 435134
rect 64258 434898 64342 435134
rect 64578 434898 64662 435134
rect 64898 434898 64982 435134
rect 65218 434898 65302 435134
rect 65538 434898 65622 435134
rect 65858 434898 65960 435134
rect 62960 434866 65960 434898
rect 71801 435454 72149 435486
rect 71801 435218 71857 435454
rect 72093 435218 72149 435454
rect 71801 435134 72149 435218
rect 71801 434898 71857 435134
rect 72093 434898 72149 435134
rect 71801 434866 72149 434898
rect 165505 435454 165853 435486
rect 165505 435218 165561 435454
rect 165797 435218 165853 435454
rect 165505 435134 165853 435218
rect 165505 434898 165561 435134
rect 165797 434898 165853 435134
rect 165505 434866 165853 434898
rect 403757 435454 404105 435486
rect 403757 435218 403813 435454
rect 404049 435218 404105 435454
rect 403757 435134 404105 435218
rect 403757 434898 403813 435134
rect 404049 434898 404105 435134
rect 403757 434866 404105 434898
rect 497461 435454 497809 435486
rect 497461 435218 497517 435454
rect 497753 435218 497809 435454
rect 497461 435134 497809 435218
rect 497461 434898 497517 435134
rect 497753 434898 497809 435134
rect 497461 434866 497809 434898
rect 503948 435454 506948 435486
rect 503948 435218 504050 435454
rect 504286 435218 504370 435454
rect 504606 435218 504690 435454
rect 504926 435218 505010 435454
rect 505246 435218 505330 435454
rect 505566 435218 505650 435454
rect 505886 435218 505970 435454
rect 506206 435218 506290 435454
rect 506526 435218 506610 435454
rect 506846 435218 506948 435454
rect 503948 435134 506948 435218
rect 503948 434898 504050 435134
rect 504286 434898 504370 435134
rect 504606 434898 504690 435134
rect 504926 434898 505010 435134
rect 505246 434898 505330 435134
rect 505566 434898 505650 435134
rect 505886 434898 505970 435134
rect 506206 434898 506290 435134
rect 506526 434898 506610 435134
rect 506846 434898 506948 435134
rect 503948 434866 506948 434898
rect 58960 417454 61960 417486
rect 58960 417218 59062 417454
rect 59298 417218 59382 417454
rect 59618 417218 59702 417454
rect 59938 417218 60022 417454
rect 60258 417218 60342 417454
rect 60578 417218 60662 417454
rect 60898 417218 60982 417454
rect 61218 417218 61302 417454
rect 61538 417218 61622 417454
rect 61858 417218 61960 417454
rect 58960 417134 61960 417218
rect 58960 416898 59062 417134
rect 59298 416898 59382 417134
rect 59618 416898 59702 417134
rect 59938 416898 60022 417134
rect 60258 416898 60342 417134
rect 60578 416898 60662 417134
rect 60898 416898 60982 417134
rect 61218 416898 61302 417134
rect 61538 416898 61622 417134
rect 61858 416898 61960 417134
rect 58960 416866 61960 416898
rect 71121 417454 71469 417486
rect 71121 417218 71177 417454
rect 71413 417218 71469 417454
rect 71121 417134 71469 417218
rect 71121 416898 71177 417134
rect 71413 416898 71469 417134
rect 71121 416866 71469 416898
rect 166185 417454 166533 417486
rect 166185 417218 166241 417454
rect 166477 417218 166533 417454
rect 166185 417134 166533 417218
rect 166185 416898 166241 417134
rect 166477 416898 166533 417134
rect 166185 416866 166533 416898
rect 403077 417454 403425 417486
rect 403077 417218 403133 417454
rect 403369 417218 403425 417454
rect 403077 417134 403425 417218
rect 403077 416898 403133 417134
rect 403369 416898 403425 417134
rect 403077 416866 403425 416898
rect 498141 417454 498489 417486
rect 498141 417218 498197 417454
rect 498433 417218 498489 417454
rect 498141 417134 498489 417218
rect 498141 416898 498197 417134
rect 498433 416898 498489 417134
rect 498141 416866 498489 416898
rect 507948 417454 510948 417486
rect 507948 417218 508050 417454
rect 508286 417218 508370 417454
rect 508606 417218 508690 417454
rect 508926 417218 509010 417454
rect 509246 417218 509330 417454
rect 509566 417218 509650 417454
rect 509886 417218 509970 417454
rect 510206 417218 510290 417454
rect 510526 417218 510610 417454
rect 510846 417218 510948 417454
rect 507948 417134 510948 417218
rect 507948 416898 508050 417134
rect 508286 416898 508370 417134
rect 508606 416898 508690 417134
rect 508926 416898 509010 417134
rect 509246 416898 509330 417134
rect 509566 416898 509650 417134
rect 509886 416898 509970 417134
rect 510206 416898 510290 417134
rect 510526 416898 510610 417134
rect 510846 416898 510948 417134
rect 507948 416866 510948 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 62960 399454 65960 399486
rect 62960 399218 63062 399454
rect 63298 399218 63382 399454
rect 63618 399218 63702 399454
rect 63938 399218 64022 399454
rect 64258 399218 64342 399454
rect 64578 399218 64662 399454
rect 64898 399218 64982 399454
rect 65218 399218 65302 399454
rect 65538 399218 65622 399454
rect 65858 399218 65960 399454
rect 62960 399134 65960 399218
rect 62960 398898 63062 399134
rect 63298 398898 63382 399134
rect 63618 398898 63702 399134
rect 63938 398898 64022 399134
rect 64258 398898 64342 399134
rect 64578 398898 64662 399134
rect 64898 398898 64982 399134
rect 65218 398898 65302 399134
rect 65538 398898 65622 399134
rect 65858 398898 65960 399134
rect 62960 398866 65960 398898
rect 71801 399454 72149 399486
rect 71801 399218 71857 399454
rect 72093 399218 72149 399454
rect 71801 399134 72149 399218
rect 71801 398898 71857 399134
rect 72093 398898 72149 399134
rect 71801 398866 72149 398898
rect 165505 399454 165853 399486
rect 165505 399218 165561 399454
rect 165797 399218 165853 399454
rect 165505 399134 165853 399218
rect 165505 398898 165561 399134
rect 165797 398898 165853 399134
rect 165505 398866 165853 398898
rect 403757 399454 404105 399486
rect 403757 399218 403813 399454
rect 404049 399218 404105 399454
rect 403757 399134 404105 399218
rect 403757 398898 403813 399134
rect 404049 398898 404105 399134
rect 403757 398866 404105 398898
rect 497461 399454 497809 399486
rect 497461 399218 497517 399454
rect 497753 399218 497809 399454
rect 497461 399134 497809 399218
rect 497461 398898 497517 399134
rect 497753 398898 497809 399134
rect 497461 398866 497809 398898
rect 503948 399454 506948 399486
rect 503948 399218 504050 399454
rect 504286 399218 504370 399454
rect 504606 399218 504690 399454
rect 504926 399218 505010 399454
rect 505246 399218 505330 399454
rect 505566 399218 505650 399454
rect 505886 399218 505970 399454
rect 506206 399218 506290 399454
rect 506526 399218 506610 399454
rect 506846 399218 506948 399454
rect 503948 399134 506948 399218
rect 503948 398898 504050 399134
rect 504286 398898 504370 399134
rect 504606 398898 504690 399134
rect 504926 398898 505010 399134
rect 505246 398898 505330 399134
rect 505566 398898 505650 399134
rect 505886 398898 505970 399134
rect 506206 398898 506290 399134
rect 506526 398898 506610 399134
rect 506846 398898 506948 399134
rect 503948 398866 506948 398898
rect 58960 381454 61960 381486
rect 58960 381218 59062 381454
rect 59298 381218 59382 381454
rect 59618 381218 59702 381454
rect 59938 381218 60022 381454
rect 60258 381218 60342 381454
rect 60578 381218 60662 381454
rect 60898 381218 60982 381454
rect 61218 381218 61302 381454
rect 61538 381218 61622 381454
rect 61858 381218 61960 381454
rect 58960 381134 61960 381218
rect 58960 380898 59062 381134
rect 59298 380898 59382 381134
rect 59618 380898 59702 381134
rect 59938 380898 60022 381134
rect 60258 380898 60342 381134
rect 60578 380898 60662 381134
rect 60898 380898 60982 381134
rect 61218 380898 61302 381134
rect 61538 380898 61622 381134
rect 61858 380898 61960 381134
rect 58960 380866 61960 380898
rect 71121 381454 71469 381486
rect 71121 381218 71177 381454
rect 71413 381218 71469 381454
rect 71121 381134 71469 381218
rect 71121 380898 71177 381134
rect 71413 380898 71469 381134
rect 71121 380866 71469 380898
rect 166185 381454 166533 381486
rect 166185 381218 166241 381454
rect 166477 381218 166533 381454
rect 166185 381134 166533 381218
rect 166185 380898 166241 381134
rect 166477 380898 166533 381134
rect 166185 380866 166533 380898
rect 403077 381454 403425 381486
rect 403077 381218 403133 381454
rect 403369 381218 403425 381454
rect 403077 381134 403425 381218
rect 403077 380898 403133 381134
rect 403369 380898 403425 381134
rect 403077 380866 403425 380898
rect 498141 381454 498489 381486
rect 498141 381218 498197 381454
rect 498433 381218 498489 381454
rect 498141 381134 498489 381218
rect 498141 380898 498197 381134
rect 498433 380898 498489 381134
rect 498141 380866 498489 380898
rect 507948 381454 510948 381486
rect 507948 381218 508050 381454
rect 508286 381218 508370 381454
rect 508606 381218 508690 381454
rect 508926 381218 509010 381454
rect 509246 381218 509330 381454
rect 509566 381218 509650 381454
rect 509886 381218 509970 381454
rect 510206 381218 510290 381454
rect 510526 381218 510610 381454
rect 510846 381218 510948 381454
rect 507948 381134 510948 381218
rect 507948 380898 508050 381134
rect 508286 380898 508370 381134
rect 508606 380898 508690 381134
rect 508926 380898 509010 381134
rect 509246 380898 509330 381134
rect 509566 380898 509650 381134
rect 509886 380898 509970 381134
rect 510206 380898 510290 381134
rect 510526 380898 510610 381134
rect 510846 380898 510948 381134
rect 507948 380866 510948 380898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 62960 363454 65960 363486
rect 62960 363218 63062 363454
rect 63298 363218 63382 363454
rect 63618 363218 63702 363454
rect 63938 363218 64022 363454
rect 64258 363218 64342 363454
rect 64578 363218 64662 363454
rect 64898 363218 64982 363454
rect 65218 363218 65302 363454
rect 65538 363218 65622 363454
rect 65858 363218 65960 363454
rect 62960 363134 65960 363218
rect 62960 362898 63062 363134
rect 63298 362898 63382 363134
rect 63618 362898 63702 363134
rect 63938 362898 64022 363134
rect 64258 362898 64342 363134
rect 64578 362898 64662 363134
rect 64898 362898 64982 363134
rect 65218 362898 65302 363134
rect 65538 362898 65622 363134
rect 65858 362898 65960 363134
rect 62960 362866 65960 362898
rect 503948 363454 506948 363486
rect 503948 363218 504050 363454
rect 504286 363218 504370 363454
rect 504606 363218 504690 363454
rect 504926 363218 505010 363454
rect 505246 363218 505330 363454
rect 505566 363218 505650 363454
rect 505886 363218 505970 363454
rect 506206 363218 506290 363454
rect 506526 363218 506610 363454
rect 506846 363218 506948 363454
rect 503948 363134 506948 363218
rect 503948 362898 504050 363134
rect 504286 362898 504370 363134
rect 504606 362898 504690 363134
rect 504926 362898 505010 363134
rect 505246 362898 505330 363134
rect 505566 362898 505650 363134
rect 505886 362898 505970 363134
rect 506206 362898 506290 363134
rect 506526 362898 506610 363134
rect 506846 362898 506948 363134
rect 503948 362866 506948 362898
rect 58960 345454 61960 345486
rect 58960 345218 59062 345454
rect 59298 345218 59382 345454
rect 59618 345218 59702 345454
rect 59938 345218 60022 345454
rect 60258 345218 60342 345454
rect 60578 345218 60662 345454
rect 60898 345218 60982 345454
rect 61218 345218 61302 345454
rect 61538 345218 61622 345454
rect 61858 345218 61960 345454
rect 58960 345134 61960 345218
rect 58960 344898 59062 345134
rect 59298 344898 59382 345134
rect 59618 344898 59702 345134
rect 59938 344898 60022 345134
rect 60258 344898 60342 345134
rect 60578 344898 60662 345134
rect 60898 344898 60982 345134
rect 61218 344898 61302 345134
rect 61538 344898 61622 345134
rect 61858 344898 61960 345134
rect 58960 344866 61960 344898
rect 71121 345454 71469 345486
rect 71121 345218 71177 345454
rect 71413 345218 71469 345454
rect 71121 345134 71469 345218
rect 71121 344898 71177 345134
rect 71413 344898 71469 345134
rect 71121 344866 71469 344898
rect 166185 345454 166533 345486
rect 166185 345218 166241 345454
rect 166477 345218 166533 345454
rect 166185 345134 166533 345218
rect 166185 344898 166241 345134
rect 166477 344898 166533 345134
rect 166185 344866 166533 344898
rect 403077 345454 403425 345486
rect 403077 345218 403133 345454
rect 403369 345218 403425 345454
rect 403077 345134 403425 345218
rect 403077 344898 403133 345134
rect 403369 344898 403425 345134
rect 403077 344866 403425 344898
rect 498141 345454 498489 345486
rect 498141 345218 498197 345454
rect 498433 345218 498489 345454
rect 498141 345134 498489 345218
rect 498141 344898 498197 345134
rect 498433 344898 498489 345134
rect 498141 344866 498489 344898
rect 507948 345454 510948 345486
rect 507948 345218 508050 345454
rect 508286 345218 508370 345454
rect 508606 345218 508690 345454
rect 508926 345218 509010 345454
rect 509246 345218 509330 345454
rect 509566 345218 509650 345454
rect 509886 345218 509970 345454
rect 510206 345218 510290 345454
rect 510526 345218 510610 345454
rect 510846 345218 510948 345454
rect 507948 345134 510948 345218
rect 507948 344898 508050 345134
rect 508286 344898 508370 345134
rect 508606 344898 508690 345134
rect 508926 344898 509010 345134
rect 509246 344898 509330 345134
rect 509566 344898 509650 345134
rect 509886 344898 509970 345134
rect 510206 344898 510290 345134
rect 510526 344898 510610 345134
rect 510846 344898 510948 345134
rect 507948 344866 510948 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 62960 327454 65960 327486
rect 62960 327218 63062 327454
rect 63298 327218 63382 327454
rect 63618 327218 63702 327454
rect 63938 327218 64022 327454
rect 64258 327218 64342 327454
rect 64578 327218 64662 327454
rect 64898 327218 64982 327454
rect 65218 327218 65302 327454
rect 65538 327218 65622 327454
rect 65858 327218 65960 327454
rect 62960 327134 65960 327218
rect 62960 326898 63062 327134
rect 63298 326898 63382 327134
rect 63618 326898 63702 327134
rect 63938 326898 64022 327134
rect 64258 326898 64342 327134
rect 64578 326898 64662 327134
rect 64898 326898 64982 327134
rect 65218 326898 65302 327134
rect 65538 326898 65622 327134
rect 65858 326898 65960 327134
rect 62960 326866 65960 326898
rect 71801 327454 72149 327486
rect 71801 327218 71857 327454
rect 72093 327218 72149 327454
rect 71801 327134 72149 327218
rect 71801 326898 71857 327134
rect 72093 326898 72149 327134
rect 71801 326866 72149 326898
rect 165505 327454 165853 327486
rect 165505 327218 165561 327454
rect 165797 327218 165853 327454
rect 165505 327134 165853 327218
rect 165505 326898 165561 327134
rect 165797 326898 165853 327134
rect 165505 326866 165853 326898
rect 403757 327454 404105 327486
rect 403757 327218 403813 327454
rect 404049 327218 404105 327454
rect 403757 327134 404105 327218
rect 403757 326898 403813 327134
rect 404049 326898 404105 327134
rect 403757 326866 404105 326898
rect 497461 327454 497809 327486
rect 497461 327218 497517 327454
rect 497753 327218 497809 327454
rect 497461 327134 497809 327218
rect 497461 326898 497517 327134
rect 497753 326898 497809 327134
rect 497461 326866 497809 326898
rect 503948 327454 506948 327486
rect 503948 327218 504050 327454
rect 504286 327218 504370 327454
rect 504606 327218 504690 327454
rect 504926 327218 505010 327454
rect 505246 327218 505330 327454
rect 505566 327218 505650 327454
rect 505886 327218 505970 327454
rect 506206 327218 506290 327454
rect 506526 327218 506610 327454
rect 506846 327218 506948 327454
rect 503948 327134 506948 327218
rect 503948 326898 504050 327134
rect 504286 326898 504370 327134
rect 504606 326898 504690 327134
rect 504926 326898 505010 327134
rect 505246 326898 505330 327134
rect 505566 326898 505650 327134
rect 505886 326898 505970 327134
rect 506206 326898 506290 327134
rect 506526 326898 506610 327134
rect 506846 326898 506948 327134
rect 503948 326866 506948 326898
rect 58960 309454 61960 309486
rect 58960 309218 59062 309454
rect 59298 309218 59382 309454
rect 59618 309218 59702 309454
rect 59938 309218 60022 309454
rect 60258 309218 60342 309454
rect 60578 309218 60662 309454
rect 60898 309218 60982 309454
rect 61218 309218 61302 309454
rect 61538 309218 61622 309454
rect 61858 309218 61960 309454
rect 58960 309134 61960 309218
rect 58960 308898 59062 309134
rect 59298 308898 59382 309134
rect 59618 308898 59702 309134
rect 59938 308898 60022 309134
rect 60258 308898 60342 309134
rect 60578 308898 60662 309134
rect 60898 308898 60982 309134
rect 61218 308898 61302 309134
rect 61538 308898 61622 309134
rect 61858 308898 61960 309134
rect 58960 308866 61960 308898
rect 71121 309454 71469 309486
rect 71121 309218 71177 309454
rect 71413 309218 71469 309454
rect 71121 309134 71469 309218
rect 71121 308898 71177 309134
rect 71413 308898 71469 309134
rect 71121 308866 71469 308898
rect 166185 309454 166533 309486
rect 166185 309218 166241 309454
rect 166477 309218 166533 309454
rect 166185 309134 166533 309218
rect 166185 308898 166241 309134
rect 166477 308898 166533 309134
rect 166185 308866 166533 308898
rect 403077 309454 403425 309486
rect 403077 309218 403133 309454
rect 403369 309218 403425 309454
rect 403077 309134 403425 309218
rect 403077 308898 403133 309134
rect 403369 308898 403425 309134
rect 403077 308866 403425 308898
rect 498141 309454 498489 309486
rect 498141 309218 498197 309454
rect 498433 309218 498489 309454
rect 498141 309134 498489 309218
rect 498141 308898 498197 309134
rect 498433 308898 498489 309134
rect 498141 308866 498489 308898
rect 507948 309454 510948 309486
rect 507948 309218 508050 309454
rect 508286 309218 508370 309454
rect 508606 309218 508690 309454
rect 508926 309218 509010 309454
rect 509246 309218 509330 309454
rect 509566 309218 509650 309454
rect 509886 309218 509970 309454
rect 510206 309218 510290 309454
rect 510526 309218 510610 309454
rect 510846 309218 510948 309454
rect 507948 309134 510948 309218
rect 507948 308898 508050 309134
rect 508286 308898 508370 309134
rect 508606 308898 508690 309134
rect 508926 308898 509010 309134
rect 509246 308898 509330 309134
rect 509566 308898 509650 309134
rect 509886 308898 509970 309134
rect 510206 308898 510290 309134
rect 510526 308898 510610 309134
rect 510846 308898 510948 309134
rect 507948 308866 510948 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 62960 291454 65960 291486
rect 62960 291218 63062 291454
rect 63298 291218 63382 291454
rect 63618 291218 63702 291454
rect 63938 291218 64022 291454
rect 64258 291218 64342 291454
rect 64578 291218 64662 291454
rect 64898 291218 64982 291454
rect 65218 291218 65302 291454
rect 65538 291218 65622 291454
rect 65858 291218 65960 291454
rect 62960 291134 65960 291218
rect 62960 290898 63062 291134
rect 63298 290898 63382 291134
rect 63618 290898 63702 291134
rect 63938 290898 64022 291134
rect 64258 290898 64342 291134
rect 64578 290898 64662 291134
rect 64898 290898 64982 291134
rect 65218 290898 65302 291134
rect 65538 290898 65622 291134
rect 65858 290898 65960 291134
rect 62960 290866 65960 290898
rect 71801 291454 72149 291486
rect 71801 291218 71857 291454
rect 72093 291218 72149 291454
rect 71801 291134 72149 291218
rect 71801 290898 71857 291134
rect 72093 290898 72149 291134
rect 71801 290866 72149 290898
rect 165505 291454 165853 291486
rect 165505 291218 165561 291454
rect 165797 291218 165853 291454
rect 165505 291134 165853 291218
rect 165505 290898 165561 291134
rect 165797 290898 165853 291134
rect 165505 290866 165853 290898
rect 403757 291454 404105 291486
rect 403757 291218 403813 291454
rect 404049 291218 404105 291454
rect 403757 291134 404105 291218
rect 403757 290898 403813 291134
rect 404049 290898 404105 291134
rect 403757 290866 404105 290898
rect 497461 291454 497809 291486
rect 497461 291218 497517 291454
rect 497753 291218 497809 291454
rect 497461 291134 497809 291218
rect 497461 290898 497517 291134
rect 497753 290898 497809 291134
rect 497461 290866 497809 290898
rect 503948 291454 506948 291486
rect 503948 291218 504050 291454
rect 504286 291218 504370 291454
rect 504606 291218 504690 291454
rect 504926 291218 505010 291454
rect 505246 291218 505330 291454
rect 505566 291218 505650 291454
rect 505886 291218 505970 291454
rect 506206 291218 506290 291454
rect 506526 291218 506610 291454
rect 506846 291218 506948 291454
rect 503948 291134 506948 291218
rect 503948 290898 504050 291134
rect 504286 290898 504370 291134
rect 504606 290898 504690 291134
rect 504926 290898 505010 291134
rect 505246 290898 505330 291134
rect 505566 290898 505650 291134
rect 505886 290898 505970 291134
rect 506206 290898 506290 291134
rect 506526 290898 506610 291134
rect 506846 290898 506948 291134
rect 503948 290866 506948 290898
rect 58960 273454 61960 273486
rect 58960 273218 59062 273454
rect 59298 273218 59382 273454
rect 59618 273218 59702 273454
rect 59938 273218 60022 273454
rect 60258 273218 60342 273454
rect 60578 273218 60662 273454
rect 60898 273218 60982 273454
rect 61218 273218 61302 273454
rect 61538 273218 61622 273454
rect 61858 273218 61960 273454
rect 58960 273134 61960 273218
rect 58960 272898 59062 273134
rect 59298 272898 59382 273134
rect 59618 272898 59702 273134
rect 59938 272898 60022 273134
rect 60258 272898 60342 273134
rect 60578 272898 60662 273134
rect 60898 272898 60982 273134
rect 61218 272898 61302 273134
rect 61538 272898 61622 273134
rect 61858 272898 61960 273134
rect 58960 272866 61960 272898
rect 507948 273454 510948 273486
rect 507948 273218 508050 273454
rect 508286 273218 508370 273454
rect 508606 273218 508690 273454
rect 508926 273218 509010 273454
rect 509246 273218 509330 273454
rect 509566 273218 509650 273454
rect 509886 273218 509970 273454
rect 510206 273218 510290 273454
rect 510526 273218 510610 273454
rect 510846 273218 510948 273454
rect 507948 273134 510948 273218
rect 507948 272898 508050 273134
rect 508286 272898 508370 273134
rect 508606 272898 508690 273134
rect 508926 272898 509010 273134
rect 509246 272898 509330 273134
rect 509566 272898 509650 273134
rect 509886 272898 509970 273134
rect 510206 272898 510290 273134
rect 510526 272898 510610 273134
rect 510846 272898 510948 273134
rect 507948 272866 510948 272898
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 62960 255454 65960 255486
rect 62960 255218 63062 255454
rect 63298 255218 63382 255454
rect 63618 255218 63702 255454
rect 63938 255218 64022 255454
rect 64258 255218 64342 255454
rect 64578 255218 64662 255454
rect 64898 255218 64982 255454
rect 65218 255218 65302 255454
rect 65538 255218 65622 255454
rect 65858 255218 65960 255454
rect 62960 255134 65960 255218
rect 62960 254898 63062 255134
rect 63298 254898 63382 255134
rect 63618 254898 63702 255134
rect 63938 254898 64022 255134
rect 64258 254898 64342 255134
rect 64578 254898 64662 255134
rect 64898 254898 64982 255134
rect 65218 254898 65302 255134
rect 65538 254898 65622 255134
rect 65858 254898 65960 255134
rect 62960 254866 65960 254898
rect 503948 255454 506948 255486
rect 503948 255218 504050 255454
rect 504286 255218 504370 255454
rect 504606 255218 504690 255454
rect 504926 255218 505010 255454
rect 505246 255218 505330 255454
rect 505566 255218 505650 255454
rect 505886 255218 505970 255454
rect 506206 255218 506290 255454
rect 506526 255218 506610 255454
rect 506846 255218 506948 255454
rect 503948 255134 506948 255218
rect 503948 254898 504050 255134
rect 504286 254898 504370 255134
rect 504606 254898 504690 255134
rect 504926 254898 505010 255134
rect 505246 254898 505330 255134
rect 505566 254898 505650 255134
rect 505886 254898 505970 255134
rect 506206 254898 506290 255134
rect 506526 254898 506610 255134
rect 506846 254898 506948 255134
rect 503948 254866 506948 254898
rect 58960 237454 61960 237486
rect 58960 237218 59062 237454
rect 59298 237218 59382 237454
rect 59618 237218 59702 237454
rect 59938 237218 60022 237454
rect 60258 237218 60342 237454
rect 60578 237218 60662 237454
rect 60898 237218 60982 237454
rect 61218 237218 61302 237454
rect 61538 237218 61622 237454
rect 61858 237218 61960 237454
rect 58960 237134 61960 237218
rect 58960 236898 59062 237134
rect 59298 236898 59382 237134
rect 59618 236898 59702 237134
rect 59938 236898 60022 237134
rect 60258 236898 60342 237134
rect 60578 236898 60662 237134
rect 60898 236898 60982 237134
rect 61218 236898 61302 237134
rect 61538 236898 61622 237134
rect 61858 236898 61960 237134
rect 58960 236866 61960 236898
rect 71121 237454 71469 237486
rect 71121 237218 71177 237454
rect 71413 237218 71469 237454
rect 71121 237134 71469 237218
rect 71121 236898 71177 237134
rect 71413 236898 71469 237134
rect 71121 236866 71469 236898
rect 166185 237454 166533 237486
rect 166185 237218 166241 237454
rect 166477 237218 166533 237454
rect 166185 237134 166533 237218
rect 166185 236898 166241 237134
rect 166477 236898 166533 237134
rect 166185 236866 166533 236898
rect 403077 237454 403425 237486
rect 403077 237218 403133 237454
rect 403369 237218 403425 237454
rect 403077 237134 403425 237218
rect 403077 236898 403133 237134
rect 403369 236898 403425 237134
rect 403077 236866 403425 236898
rect 498141 237454 498489 237486
rect 498141 237218 498197 237454
rect 498433 237218 498489 237454
rect 498141 237134 498489 237218
rect 498141 236898 498197 237134
rect 498433 236898 498489 237134
rect 498141 236866 498489 236898
rect 507948 237454 510948 237486
rect 507948 237218 508050 237454
rect 508286 237218 508370 237454
rect 508606 237218 508690 237454
rect 508926 237218 509010 237454
rect 509246 237218 509330 237454
rect 509566 237218 509650 237454
rect 509886 237218 509970 237454
rect 510206 237218 510290 237454
rect 510526 237218 510610 237454
rect 510846 237218 510948 237454
rect 507948 237134 510948 237218
rect 507948 236898 508050 237134
rect 508286 236898 508370 237134
rect 508606 236898 508690 237134
rect 508926 236898 509010 237134
rect 509246 236898 509330 237134
rect 509566 236898 509650 237134
rect 509886 236898 509970 237134
rect 510206 236898 510290 237134
rect 510526 236898 510610 237134
rect 510846 236898 510948 237134
rect 507948 236866 510948 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 62960 219454 65960 219486
rect 62960 219218 63062 219454
rect 63298 219218 63382 219454
rect 63618 219218 63702 219454
rect 63938 219218 64022 219454
rect 64258 219218 64342 219454
rect 64578 219218 64662 219454
rect 64898 219218 64982 219454
rect 65218 219218 65302 219454
rect 65538 219218 65622 219454
rect 65858 219218 65960 219454
rect 62960 219134 65960 219218
rect 62960 218898 63062 219134
rect 63298 218898 63382 219134
rect 63618 218898 63702 219134
rect 63938 218898 64022 219134
rect 64258 218898 64342 219134
rect 64578 218898 64662 219134
rect 64898 218898 64982 219134
rect 65218 218898 65302 219134
rect 65538 218898 65622 219134
rect 65858 218898 65960 219134
rect 62960 218866 65960 218898
rect 71801 219454 72149 219486
rect 71801 219218 71857 219454
rect 72093 219218 72149 219454
rect 71801 219134 72149 219218
rect 71801 218898 71857 219134
rect 72093 218898 72149 219134
rect 71801 218866 72149 218898
rect 165505 219454 165853 219486
rect 165505 219218 165561 219454
rect 165797 219218 165853 219454
rect 165505 219134 165853 219218
rect 165505 218898 165561 219134
rect 165797 218898 165853 219134
rect 165505 218866 165853 218898
rect 403757 219454 404105 219486
rect 403757 219218 403813 219454
rect 404049 219218 404105 219454
rect 403757 219134 404105 219218
rect 403757 218898 403813 219134
rect 404049 218898 404105 219134
rect 403757 218866 404105 218898
rect 497461 219454 497809 219486
rect 497461 219218 497517 219454
rect 497753 219218 497809 219454
rect 497461 219134 497809 219218
rect 497461 218898 497517 219134
rect 497753 218898 497809 219134
rect 497461 218866 497809 218898
rect 503948 219454 506948 219486
rect 503948 219218 504050 219454
rect 504286 219218 504370 219454
rect 504606 219218 504690 219454
rect 504926 219218 505010 219454
rect 505246 219218 505330 219454
rect 505566 219218 505650 219454
rect 505886 219218 505970 219454
rect 506206 219218 506290 219454
rect 506526 219218 506610 219454
rect 506846 219218 506948 219454
rect 503948 219134 506948 219218
rect 503948 218898 504050 219134
rect 504286 218898 504370 219134
rect 504606 218898 504690 219134
rect 504926 218898 505010 219134
rect 505246 218898 505330 219134
rect 505566 218898 505650 219134
rect 505886 218898 505970 219134
rect 506206 218898 506290 219134
rect 506526 218898 506610 219134
rect 506846 218898 506948 219134
rect 503948 218866 506948 218898
rect 58960 201454 61960 201486
rect 58960 201218 59062 201454
rect 59298 201218 59382 201454
rect 59618 201218 59702 201454
rect 59938 201218 60022 201454
rect 60258 201218 60342 201454
rect 60578 201218 60662 201454
rect 60898 201218 60982 201454
rect 61218 201218 61302 201454
rect 61538 201218 61622 201454
rect 61858 201218 61960 201454
rect 58960 201134 61960 201218
rect 58960 200898 59062 201134
rect 59298 200898 59382 201134
rect 59618 200898 59702 201134
rect 59938 200898 60022 201134
rect 60258 200898 60342 201134
rect 60578 200898 60662 201134
rect 60898 200898 60982 201134
rect 61218 200898 61302 201134
rect 61538 200898 61622 201134
rect 61858 200898 61960 201134
rect 58960 200866 61960 200898
rect 71121 201454 71469 201486
rect 71121 201218 71177 201454
rect 71413 201218 71469 201454
rect 71121 201134 71469 201218
rect 71121 200898 71177 201134
rect 71413 200898 71469 201134
rect 71121 200866 71469 200898
rect 166185 201454 166533 201486
rect 166185 201218 166241 201454
rect 166477 201218 166533 201454
rect 166185 201134 166533 201218
rect 166185 200898 166241 201134
rect 166477 200898 166533 201134
rect 166185 200866 166533 200898
rect 403077 201454 403425 201486
rect 403077 201218 403133 201454
rect 403369 201218 403425 201454
rect 403077 201134 403425 201218
rect 403077 200898 403133 201134
rect 403369 200898 403425 201134
rect 403077 200866 403425 200898
rect 498141 201454 498489 201486
rect 498141 201218 498197 201454
rect 498433 201218 498489 201454
rect 498141 201134 498489 201218
rect 498141 200898 498197 201134
rect 498433 200898 498489 201134
rect 498141 200866 498489 200898
rect 507948 201454 510948 201486
rect 507948 201218 508050 201454
rect 508286 201218 508370 201454
rect 508606 201218 508690 201454
rect 508926 201218 509010 201454
rect 509246 201218 509330 201454
rect 509566 201218 509650 201454
rect 509886 201218 509970 201454
rect 510206 201218 510290 201454
rect 510526 201218 510610 201454
rect 510846 201218 510948 201454
rect 507948 201134 510948 201218
rect 507948 200898 508050 201134
rect 508286 200898 508370 201134
rect 508606 200898 508690 201134
rect 508926 200898 509010 201134
rect 509246 200898 509330 201134
rect 509566 200898 509650 201134
rect 509886 200898 509970 201134
rect 510206 200898 510290 201134
rect 510526 200898 510610 201134
rect 510846 200898 510948 201134
rect 507948 200866 510948 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 62960 183454 65960 183486
rect 62960 183218 63062 183454
rect 63298 183218 63382 183454
rect 63618 183218 63702 183454
rect 63938 183218 64022 183454
rect 64258 183218 64342 183454
rect 64578 183218 64662 183454
rect 64898 183218 64982 183454
rect 65218 183218 65302 183454
rect 65538 183218 65622 183454
rect 65858 183218 65960 183454
rect 62960 183134 65960 183218
rect 62960 182898 63062 183134
rect 63298 182898 63382 183134
rect 63618 182898 63702 183134
rect 63938 182898 64022 183134
rect 64258 182898 64342 183134
rect 64578 182898 64662 183134
rect 64898 182898 64982 183134
rect 65218 182898 65302 183134
rect 65538 182898 65622 183134
rect 65858 182898 65960 183134
rect 62960 182866 65960 182898
rect 71801 183454 72149 183486
rect 71801 183218 71857 183454
rect 72093 183218 72149 183454
rect 71801 183134 72149 183218
rect 71801 182898 71857 183134
rect 72093 182898 72149 183134
rect 71801 182866 72149 182898
rect 165505 183454 165853 183486
rect 165505 183218 165561 183454
rect 165797 183218 165853 183454
rect 165505 183134 165853 183218
rect 165505 182898 165561 183134
rect 165797 182898 165853 183134
rect 165505 182866 165853 182898
rect 403757 183454 404105 183486
rect 403757 183218 403813 183454
rect 404049 183218 404105 183454
rect 403757 183134 404105 183218
rect 403757 182898 403813 183134
rect 404049 182898 404105 183134
rect 403757 182866 404105 182898
rect 497461 183454 497809 183486
rect 497461 183218 497517 183454
rect 497753 183218 497809 183454
rect 497461 183134 497809 183218
rect 497461 182898 497517 183134
rect 497753 182898 497809 183134
rect 497461 182866 497809 182898
rect 503948 183454 506948 183486
rect 503948 183218 504050 183454
rect 504286 183218 504370 183454
rect 504606 183218 504690 183454
rect 504926 183218 505010 183454
rect 505246 183218 505330 183454
rect 505566 183218 505650 183454
rect 505886 183218 505970 183454
rect 506206 183218 506290 183454
rect 506526 183218 506610 183454
rect 506846 183218 506948 183454
rect 503948 183134 506948 183218
rect 503948 182898 504050 183134
rect 504286 182898 504370 183134
rect 504606 182898 504690 183134
rect 504926 182898 505010 183134
rect 505246 182898 505330 183134
rect 505566 182898 505650 183134
rect 505886 182898 505970 183134
rect 506206 182898 506290 183134
rect 506526 182898 506610 183134
rect 506846 182898 506948 183134
rect 503948 182866 506948 182898
rect 58960 165454 61960 165486
rect 58960 165218 59062 165454
rect 59298 165218 59382 165454
rect 59618 165218 59702 165454
rect 59938 165218 60022 165454
rect 60258 165218 60342 165454
rect 60578 165218 60662 165454
rect 60898 165218 60982 165454
rect 61218 165218 61302 165454
rect 61538 165218 61622 165454
rect 61858 165218 61960 165454
rect 58960 165134 61960 165218
rect 58960 164898 59062 165134
rect 59298 164898 59382 165134
rect 59618 164898 59702 165134
rect 59938 164898 60022 165134
rect 60258 164898 60342 165134
rect 60578 164898 60662 165134
rect 60898 164898 60982 165134
rect 61218 164898 61302 165134
rect 61538 164898 61622 165134
rect 61858 164898 61960 165134
rect 58960 164866 61960 164898
rect 507948 165454 510948 165486
rect 507948 165218 508050 165454
rect 508286 165218 508370 165454
rect 508606 165218 508690 165454
rect 508926 165218 509010 165454
rect 509246 165218 509330 165454
rect 509566 165218 509650 165454
rect 509886 165218 509970 165454
rect 510206 165218 510290 165454
rect 510526 165218 510610 165454
rect 510846 165218 510948 165454
rect 507948 165134 510948 165218
rect 507948 164898 508050 165134
rect 508286 164898 508370 165134
rect 508606 164898 508690 165134
rect 508926 164898 509010 165134
rect 509246 164898 509330 165134
rect 509566 164898 509650 165134
rect 509886 164898 509970 165134
rect 510206 164898 510290 165134
rect 510526 164898 510610 165134
rect 510846 164898 510948 165134
rect 507948 164866 510948 164898
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 62960 147454 65960 147486
rect 62960 147218 63062 147454
rect 63298 147218 63382 147454
rect 63618 147218 63702 147454
rect 63938 147218 64022 147454
rect 64258 147218 64342 147454
rect 64578 147218 64662 147454
rect 64898 147218 64982 147454
rect 65218 147218 65302 147454
rect 65538 147218 65622 147454
rect 65858 147218 65960 147454
rect 62960 147134 65960 147218
rect 62960 146898 63062 147134
rect 63298 146898 63382 147134
rect 63618 146898 63702 147134
rect 63938 146898 64022 147134
rect 64258 146898 64342 147134
rect 64578 146898 64662 147134
rect 64898 146898 64982 147134
rect 65218 146898 65302 147134
rect 65538 146898 65622 147134
rect 65858 146898 65960 147134
rect 62960 146866 65960 146898
rect 71801 147454 72149 147486
rect 71801 147218 71857 147454
rect 72093 147218 72149 147454
rect 71801 147134 72149 147218
rect 71801 146898 71857 147134
rect 72093 146898 72149 147134
rect 71801 146866 72149 146898
rect 165505 147454 165853 147486
rect 165505 147218 165561 147454
rect 165797 147218 165853 147454
rect 165505 147134 165853 147218
rect 165505 146898 165561 147134
rect 165797 146898 165853 147134
rect 165505 146866 165853 146898
rect 403757 147454 404105 147486
rect 403757 147218 403813 147454
rect 404049 147218 404105 147454
rect 403757 147134 404105 147218
rect 403757 146898 403813 147134
rect 404049 146898 404105 147134
rect 403757 146866 404105 146898
rect 497461 147454 497809 147486
rect 497461 147218 497517 147454
rect 497753 147218 497809 147454
rect 497461 147134 497809 147218
rect 497461 146898 497517 147134
rect 497753 146898 497809 147134
rect 497461 146866 497809 146898
rect 503948 147454 506948 147486
rect 503948 147218 504050 147454
rect 504286 147218 504370 147454
rect 504606 147218 504690 147454
rect 504926 147218 505010 147454
rect 505246 147218 505330 147454
rect 505566 147218 505650 147454
rect 505886 147218 505970 147454
rect 506206 147218 506290 147454
rect 506526 147218 506610 147454
rect 506846 147218 506948 147454
rect 503948 147134 506948 147218
rect 503948 146898 504050 147134
rect 504286 146898 504370 147134
rect 504606 146898 504690 147134
rect 504926 146898 505010 147134
rect 505246 146898 505330 147134
rect 505566 146898 505650 147134
rect 505886 146898 505970 147134
rect 506206 146898 506290 147134
rect 506526 146898 506610 147134
rect 506846 146898 506948 147134
rect 503948 146866 506948 146898
rect 58960 129454 61960 129486
rect 58960 129218 59062 129454
rect 59298 129218 59382 129454
rect 59618 129218 59702 129454
rect 59938 129218 60022 129454
rect 60258 129218 60342 129454
rect 60578 129218 60662 129454
rect 60898 129218 60982 129454
rect 61218 129218 61302 129454
rect 61538 129218 61622 129454
rect 61858 129218 61960 129454
rect 58960 129134 61960 129218
rect 58960 128898 59062 129134
rect 59298 128898 59382 129134
rect 59618 128898 59702 129134
rect 59938 128898 60022 129134
rect 60258 128898 60342 129134
rect 60578 128898 60662 129134
rect 60898 128898 60982 129134
rect 61218 128898 61302 129134
rect 61538 128898 61622 129134
rect 61858 128898 61960 129134
rect 58960 128866 61960 128898
rect 71121 129454 71469 129486
rect 71121 129218 71177 129454
rect 71413 129218 71469 129454
rect 71121 129134 71469 129218
rect 71121 128898 71177 129134
rect 71413 128898 71469 129134
rect 71121 128866 71469 128898
rect 166185 129454 166533 129486
rect 166185 129218 166241 129454
rect 166477 129218 166533 129454
rect 166185 129134 166533 129218
rect 166185 128898 166241 129134
rect 166477 128898 166533 129134
rect 166185 128866 166533 128898
rect 403077 129454 403425 129486
rect 403077 129218 403133 129454
rect 403369 129218 403425 129454
rect 403077 129134 403425 129218
rect 403077 128898 403133 129134
rect 403369 128898 403425 129134
rect 403077 128866 403425 128898
rect 498141 129454 498489 129486
rect 498141 129218 498197 129454
rect 498433 129218 498489 129454
rect 498141 129134 498489 129218
rect 498141 128898 498197 129134
rect 498433 128898 498489 129134
rect 498141 128866 498489 128898
rect 507948 129454 510948 129486
rect 507948 129218 508050 129454
rect 508286 129218 508370 129454
rect 508606 129218 508690 129454
rect 508926 129218 509010 129454
rect 509246 129218 509330 129454
rect 509566 129218 509650 129454
rect 509886 129218 509970 129454
rect 510206 129218 510290 129454
rect 510526 129218 510610 129454
rect 510846 129218 510948 129454
rect 507948 129134 510948 129218
rect 507948 128898 508050 129134
rect 508286 128898 508370 129134
rect 508606 128898 508690 129134
rect 508926 128898 509010 129134
rect 509246 128898 509330 129134
rect 509566 128898 509650 129134
rect 509886 128898 509970 129134
rect 510206 128898 510290 129134
rect 510526 128898 510610 129134
rect 510846 128898 510948 129134
rect 507948 128866 510948 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 62960 111454 65960 111486
rect 62960 111218 63062 111454
rect 63298 111218 63382 111454
rect 63618 111218 63702 111454
rect 63938 111218 64022 111454
rect 64258 111218 64342 111454
rect 64578 111218 64662 111454
rect 64898 111218 64982 111454
rect 65218 111218 65302 111454
rect 65538 111218 65622 111454
rect 65858 111218 65960 111454
rect 62960 111134 65960 111218
rect 62960 110898 63062 111134
rect 63298 110898 63382 111134
rect 63618 110898 63702 111134
rect 63938 110898 64022 111134
rect 64258 110898 64342 111134
rect 64578 110898 64662 111134
rect 64898 110898 64982 111134
rect 65218 110898 65302 111134
rect 65538 110898 65622 111134
rect 65858 110898 65960 111134
rect 62960 110866 65960 110898
rect 71801 111454 72149 111486
rect 71801 111218 71857 111454
rect 72093 111218 72149 111454
rect 71801 111134 72149 111218
rect 71801 110898 71857 111134
rect 72093 110898 72149 111134
rect 71801 110866 72149 110898
rect 165505 111454 165853 111486
rect 165505 111218 165561 111454
rect 165797 111218 165853 111454
rect 165505 111134 165853 111218
rect 165505 110898 165561 111134
rect 165797 110898 165853 111134
rect 165505 110866 165853 110898
rect 403757 111454 404105 111486
rect 403757 111218 403813 111454
rect 404049 111218 404105 111454
rect 403757 111134 404105 111218
rect 403757 110898 403813 111134
rect 404049 110898 404105 111134
rect 403757 110866 404105 110898
rect 497461 111454 497809 111486
rect 497461 111218 497517 111454
rect 497753 111218 497809 111454
rect 497461 111134 497809 111218
rect 497461 110898 497517 111134
rect 497753 110898 497809 111134
rect 497461 110866 497809 110898
rect 503948 111454 506948 111486
rect 503948 111218 504050 111454
rect 504286 111218 504370 111454
rect 504606 111218 504690 111454
rect 504926 111218 505010 111454
rect 505246 111218 505330 111454
rect 505566 111218 505650 111454
rect 505886 111218 505970 111454
rect 506206 111218 506290 111454
rect 506526 111218 506610 111454
rect 506846 111218 506948 111454
rect 503948 111134 506948 111218
rect 503948 110898 504050 111134
rect 504286 110898 504370 111134
rect 504606 110898 504690 111134
rect 504926 110898 505010 111134
rect 505246 110898 505330 111134
rect 505566 110898 505650 111134
rect 505886 110898 505970 111134
rect 506206 110898 506290 111134
rect 506526 110898 506610 111134
rect 506846 110898 506948 111134
rect 503948 110866 506948 110898
rect 58960 93454 61960 93486
rect 58960 93218 59062 93454
rect 59298 93218 59382 93454
rect 59618 93218 59702 93454
rect 59938 93218 60022 93454
rect 60258 93218 60342 93454
rect 60578 93218 60662 93454
rect 60898 93218 60982 93454
rect 61218 93218 61302 93454
rect 61538 93218 61622 93454
rect 61858 93218 61960 93454
rect 58960 93134 61960 93218
rect 58960 92898 59062 93134
rect 59298 92898 59382 93134
rect 59618 92898 59702 93134
rect 59938 92898 60022 93134
rect 60258 92898 60342 93134
rect 60578 92898 60662 93134
rect 60898 92898 60982 93134
rect 61218 92898 61302 93134
rect 61538 92898 61622 93134
rect 61858 92898 61960 93134
rect 58960 92866 61960 92898
rect 71121 93454 71469 93486
rect 71121 93218 71177 93454
rect 71413 93218 71469 93454
rect 71121 93134 71469 93218
rect 71121 92898 71177 93134
rect 71413 92898 71469 93134
rect 71121 92866 71469 92898
rect 166185 93454 166533 93486
rect 166185 93218 166241 93454
rect 166477 93218 166533 93454
rect 166185 93134 166533 93218
rect 166185 92898 166241 93134
rect 166477 92898 166533 93134
rect 166185 92866 166533 92898
rect 403077 93454 403425 93486
rect 403077 93218 403133 93454
rect 403369 93218 403425 93454
rect 403077 93134 403425 93218
rect 403077 92898 403133 93134
rect 403369 92898 403425 93134
rect 403077 92866 403425 92898
rect 498141 93454 498489 93486
rect 498141 93218 498197 93454
rect 498433 93218 498489 93454
rect 498141 93134 498489 93218
rect 498141 92898 498197 93134
rect 498433 92898 498489 93134
rect 498141 92866 498489 92898
rect 507948 93454 510948 93486
rect 507948 93218 508050 93454
rect 508286 93218 508370 93454
rect 508606 93218 508690 93454
rect 508926 93218 509010 93454
rect 509246 93218 509330 93454
rect 509566 93218 509650 93454
rect 509886 93218 509970 93454
rect 510206 93218 510290 93454
rect 510526 93218 510610 93454
rect 510846 93218 510948 93454
rect 507948 93134 510948 93218
rect 507948 92898 508050 93134
rect 508286 92898 508370 93134
rect 508606 92898 508690 93134
rect 508926 92898 509010 93134
rect 509246 92898 509330 93134
rect 509566 92898 509650 93134
rect 509886 92898 509970 93134
rect 510206 92898 510290 93134
rect 510526 92898 510610 93134
rect 510846 92898 510948 93134
rect 507948 92866 510948 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 62960 75454 65960 75486
rect 62960 75218 63062 75454
rect 63298 75218 63382 75454
rect 63618 75218 63702 75454
rect 63938 75218 64022 75454
rect 64258 75218 64342 75454
rect 64578 75218 64662 75454
rect 64898 75218 64982 75454
rect 65218 75218 65302 75454
rect 65538 75218 65622 75454
rect 65858 75218 65960 75454
rect 62960 75134 65960 75218
rect 62960 74898 63062 75134
rect 63298 74898 63382 75134
rect 63618 74898 63702 75134
rect 63938 74898 64022 75134
rect 64258 74898 64342 75134
rect 64578 74898 64662 75134
rect 64898 74898 64982 75134
rect 65218 74898 65302 75134
rect 65538 74898 65622 75134
rect 65858 74898 65960 75134
rect 62960 74866 65960 74898
rect 503948 75454 506948 75486
rect 503948 75218 504050 75454
rect 504286 75218 504370 75454
rect 504606 75218 504690 75454
rect 504926 75218 505010 75454
rect 505246 75218 505330 75454
rect 505566 75218 505650 75454
rect 505886 75218 505970 75454
rect 506206 75218 506290 75454
rect 506526 75218 506610 75454
rect 506846 75218 506948 75454
rect 503948 75134 506948 75218
rect 503948 74898 504050 75134
rect 504286 74898 504370 75134
rect 504606 74898 504690 75134
rect 504926 74898 505010 75134
rect 505246 74898 505330 75134
rect 505566 74898 505650 75134
rect 505886 74898 505970 75134
rect 506206 74898 506290 75134
rect 506526 74898 506610 75134
rect 506846 74898 506948 75134
rect 503948 74866 506948 74898
rect 58960 57454 61960 57486
rect 58960 57218 59062 57454
rect 59298 57218 59382 57454
rect 59618 57218 59702 57454
rect 59938 57218 60022 57454
rect 60258 57218 60342 57454
rect 60578 57218 60662 57454
rect 60898 57218 60982 57454
rect 61218 57218 61302 57454
rect 61538 57218 61622 57454
rect 61858 57218 61960 57454
rect 58960 57134 61960 57218
rect 58960 56898 59062 57134
rect 59298 56898 59382 57134
rect 59618 56898 59702 57134
rect 59938 56898 60022 57134
rect 60258 56898 60342 57134
rect 60578 56898 60662 57134
rect 60898 56898 60982 57134
rect 61218 56898 61302 57134
rect 61538 56898 61622 57134
rect 61858 56898 61960 57134
rect 58960 56866 61960 56898
rect 507948 57454 510948 57486
rect 507948 57218 508050 57454
rect 508286 57218 508370 57454
rect 508606 57218 508690 57454
rect 508926 57218 509010 57454
rect 509246 57218 509330 57454
rect 509566 57218 509650 57454
rect 509886 57218 509970 57454
rect 510206 57218 510290 57454
rect 510526 57218 510610 57454
rect 510846 57218 510948 57454
rect 507948 57134 510948 57218
rect 507948 56898 508050 57134
rect 508286 56898 508370 57134
rect 508606 56898 508690 57134
rect 508926 56898 509010 57134
rect 509246 56898 509330 57134
rect 509566 56898 509650 57134
rect 509886 56898 509970 57134
rect 510206 56898 510290 57134
rect 510526 56898 510610 57134
rect 510846 56898 510948 57134
rect 507948 56866 510948 56898
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 62960 39454 65960 39486
rect 62960 39218 63062 39454
rect 63298 39218 63382 39454
rect 63618 39218 63702 39454
rect 63938 39218 64022 39454
rect 64258 39218 64342 39454
rect 64578 39218 64662 39454
rect 64898 39218 64982 39454
rect 65218 39218 65302 39454
rect 65538 39218 65622 39454
rect 65858 39218 65960 39454
rect 62960 39134 65960 39218
rect 62960 38898 63062 39134
rect 63298 38898 63382 39134
rect 63618 38898 63702 39134
rect 63938 38898 64022 39134
rect 64258 38898 64342 39134
rect 64578 38898 64662 39134
rect 64898 38898 64982 39134
rect 65218 38898 65302 39134
rect 65538 38898 65622 39134
rect 65858 38898 65960 39134
rect 62960 38866 65960 38898
rect 503948 39454 506948 39486
rect 503948 39218 504050 39454
rect 504286 39218 504370 39454
rect 504606 39218 504690 39454
rect 504926 39218 505010 39454
rect 505246 39218 505330 39454
rect 505566 39218 505650 39454
rect 505886 39218 505970 39454
rect 506206 39218 506290 39454
rect 506526 39218 506610 39454
rect 506846 39218 506948 39454
rect 503948 39134 506948 39218
rect 503948 38898 504050 39134
rect 504286 38898 504370 39134
rect 504606 38898 504690 39134
rect 504926 38898 505010 39134
rect 505246 38898 505330 39134
rect 505566 38898 505650 39134
rect 505886 38898 505970 39134
rect 506206 38898 506290 39134
rect 506526 38898 506610 39134
rect 506846 38898 506948 39134
rect 503948 38866 506948 38898
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 28000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 28000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 28000
rect 73794 3454 74414 28000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 28000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 28000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 28000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 28000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 28000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 28000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 28000
rect 109794 3454 110414 28000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 28000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 28000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 28000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 28000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 28000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 28000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 28000
rect 145794 3454 146414 28000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 28000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 28000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 28000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 28000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 28000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 28000
rect 181794 3454 182414 28000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 28000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 28000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 28000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 28000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 28000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 28000
rect 217794 3454 218414 28000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 28000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 28000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 28000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 28000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 28000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 28000
rect 253794 3454 254414 28000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 28000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 28000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 28000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 28000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 28000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 28000
rect 289794 3454 290414 28000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 28000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 28000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 28000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 28000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 28000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 28000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 28000
rect 325794 3454 326414 28000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 28000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 28000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 28000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 28000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 28000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 28000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 28000
rect 361794 3454 362414 28000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 28000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 28000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 28000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 28000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 28000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 28000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 28000
rect 397794 3454 398414 28000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 28000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 28000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 28000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 28000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 28000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 28000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 28000
rect 433794 3454 434414 28000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 28000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 28000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 28000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 28000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 28000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 28000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 28000
rect 469794 3454 470414 28000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 28000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 28000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 28000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 28000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 28000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 28000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 28000
rect 505794 3454 506414 28000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 28000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 28000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 28000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 59062 453218 59298 453454
rect 59382 453218 59618 453454
rect 59702 453218 59938 453454
rect 60022 453218 60258 453454
rect 60342 453218 60578 453454
rect 60662 453218 60898 453454
rect 60982 453218 61218 453454
rect 61302 453218 61538 453454
rect 61622 453218 61858 453454
rect 59062 452898 59298 453134
rect 59382 452898 59618 453134
rect 59702 452898 59938 453134
rect 60022 452898 60258 453134
rect 60342 452898 60578 453134
rect 60662 452898 60898 453134
rect 60982 452898 61218 453134
rect 61302 452898 61538 453134
rect 61622 452898 61858 453134
rect 71177 453218 71413 453454
rect 71177 452898 71413 453134
rect 166241 453218 166477 453454
rect 166241 452898 166477 453134
rect 403133 453218 403369 453454
rect 403133 452898 403369 453134
rect 498197 453218 498433 453454
rect 498197 452898 498433 453134
rect 508050 453218 508286 453454
rect 508370 453218 508606 453454
rect 508690 453218 508926 453454
rect 509010 453218 509246 453454
rect 509330 453218 509566 453454
rect 509650 453218 509886 453454
rect 509970 453218 510206 453454
rect 510290 453218 510526 453454
rect 510610 453218 510846 453454
rect 508050 452898 508286 453134
rect 508370 452898 508606 453134
rect 508690 452898 508926 453134
rect 509010 452898 509246 453134
rect 509330 452898 509566 453134
rect 509650 452898 509886 453134
rect 509970 452898 510206 453134
rect 510290 452898 510526 453134
rect 510610 452898 510846 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 63062 435218 63298 435454
rect 63382 435218 63618 435454
rect 63702 435218 63938 435454
rect 64022 435218 64258 435454
rect 64342 435218 64578 435454
rect 64662 435218 64898 435454
rect 64982 435218 65218 435454
rect 65302 435218 65538 435454
rect 65622 435218 65858 435454
rect 63062 434898 63298 435134
rect 63382 434898 63618 435134
rect 63702 434898 63938 435134
rect 64022 434898 64258 435134
rect 64342 434898 64578 435134
rect 64662 434898 64898 435134
rect 64982 434898 65218 435134
rect 65302 434898 65538 435134
rect 65622 434898 65858 435134
rect 71857 435218 72093 435454
rect 71857 434898 72093 435134
rect 165561 435218 165797 435454
rect 165561 434898 165797 435134
rect 403813 435218 404049 435454
rect 403813 434898 404049 435134
rect 497517 435218 497753 435454
rect 497517 434898 497753 435134
rect 504050 435218 504286 435454
rect 504370 435218 504606 435454
rect 504690 435218 504926 435454
rect 505010 435218 505246 435454
rect 505330 435218 505566 435454
rect 505650 435218 505886 435454
rect 505970 435218 506206 435454
rect 506290 435218 506526 435454
rect 506610 435218 506846 435454
rect 504050 434898 504286 435134
rect 504370 434898 504606 435134
rect 504690 434898 504926 435134
rect 505010 434898 505246 435134
rect 505330 434898 505566 435134
rect 505650 434898 505886 435134
rect 505970 434898 506206 435134
rect 506290 434898 506526 435134
rect 506610 434898 506846 435134
rect 59062 417218 59298 417454
rect 59382 417218 59618 417454
rect 59702 417218 59938 417454
rect 60022 417218 60258 417454
rect 60342 417218 60578 417454
rect 60662 417218 60898 417454
rect 60982 417218 61218 417454
rect 61302 417218 61538 417454
rect 61622 417218 61858 417454
rect 59062 416898 59298 417134
rect 59382 416898 59618 417134
rect 59702 416898 59938 417134
rect 60022 416898 60258 417134
rect 60342 416898 60578 417134
rect 60662 416898 60898 417134
rect 60982 416898 61218 417134
rect 61302 416898 61538 417134
rect 61622 416898 61858 417134
rect 71177 417218 71413 417454
rect 71177 416898 71413 417134
rect 166241 417218 166477 417454
rect 166241 416898 166477 417134
rect 403133 417218 403369 417454
rect 403133 416898 403369 417134
rect 498197 417218 498433 417454
rect 498197 416898 498433 417134
rect 508050 417218 508286 417454
rect 508370 417218 508606 417454
rect 508690 417218 508926 417454
rect 509010 417218 509246 417454
rect 509330 417218 509566 417454
rect 509650 417218 509886 417454
rect 509970 417218 510206 417454
rect 510290 417218 510526 417454
rect 510610 417218 510846 417454
rect 508050 416898 508286 417134
rect 508370 416898 508606 417134
rect 508690 416898 508926 417134
rect 509010 416898 509246 417134
rect 509330 416898 509566 417134
rect 509650 416898 509886 417134
rect 509970 416898 510206 417134
rect 510290 416898 510526 417134
rect 510610 416898 510846 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 63062 399218 63298 399454
rect 63382 399218 63618 399454
rect 63702 399218 63938 399454
rect 64022 399218 64258 399454
rect 64342 399218 64578 399454
rect 64662 399218 64898 399454
rect 64982 399218 65218 399454
rect 65302 399218 65538 399454
rect 65622 399218 65858 399454
rect 63062 398898 63298 399134
rect 63382 398898 63618 399134
rect 63702 398898 63938 399134
rect 64022 398898 64258 399134
rect 64342 398898 64578 399134
rect 64662 398898 64898 399134
rect 64982 398898 65218 399134
rect 65302 398898 65538 399134
rect 65622 398898 65858 399134
rect 71857 399218 72093 399454
rect 71857 398898 72093 399134
rect 165561 399218 165797 399454
rect 165561 398898 165797 399134
rect 403813 399218 404049 399454
rect 403813 398898 404049 399134
rect 497517 399218 497753 399454
rect 497517 398898 497753 399134
rect 504050 399218 504286 399454
rect 504370 399218 504606 399454
rect 504690 399218 504926 399454
rect 505010 399218 505246 399454
rect 505330 399218 505566 399454
rect 505650 399218 505886 399454
rect 505970 399218 506206 399454
rect 506290 399218 506526 399454
rect 506610 399218 506846 399454
rect 504050 398898 504286 399134
rect 504370 398898 504606 399134
rect 504690 398898 504926 399134
rect 505010 398898 505246 399134
rect 505330 398898 505566 399134
rect 505650 398898 505886 399134
rect 505970 398898 506206 399134
rect 506290 398898 506526 399134
rect 506610 398898 506846 399134
rect 59062 381218 59298 381454
rect 59382 381218 59618 381454
rect 59702 381218 59938 381454
rect 60022 381218 60258 381454
rect 60342 381218 60578 381454
rect 60662 381218 60898 381454
rect 60982 381218 61218 381454
rect 61302 381218 61538 381454
rect 61622 381218 61858 381454
rect 59062 380898 59298 381134
rect 59382 380898 59618 381134
rect 59702 380898 59938 381134
rect 60022 380898 60258 381134
rect 60342 380898 60578 381134
rect 60662 380898 60898 381134
rect 60982 380898 61218 381134
rect 61302 380898 61538 381134
rect 61622 380898 61858 381134
rect 71177 381218 71413 381454
rect 71177 380898 71413 381134
rect 166241 381218 166477 381454
rect 166241 380898 166477 381134
rect 403133 381218 403369 381454
rect 403133 380898 403369 381134
rect 498197 381218 498433 381454
rect 498197 380898 498433 381134
rect 508050 381218 508286 381454
rect 508370 381218 508606 381454
rect 508690 381218 508926 381454
rect 509010 381218 509246 381454
rect 509330 381218 509566 381454
rect 509650 381218 509886 381454
rect 509970 381218 510206 381454
rect 510290 381218 510526 381454
rect 510610 381218 510846 381454
rect 508050 380898 508286 381134
rect 508370 380898 508606 381134
rect 508690 380898 508926 381134
rect 509010 380898 509246 381134
rect 509330 380898 509566 381134
rect 509650 380898 509886 381134
rect 509970 380898 510206 381134
rect 510290 380898 510526 381134
rect 510610 380898 510846 381134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 63062 363218 63298 363454
rect 63382 363218 63618 363454
rect 63702 363218 63938 363454
rect 64022 363218 64258 363454
rect 64342 363218 64578 363454
rect 64662 363218 64898 363454
rect 64982 363218 65218 363454
rect 65302 363218 65538 363454
rect 65622 363218 65858 363454
rect 63062 362898 63298 363134
rect 63382 362898 63618 363134
rect 63702 362898 63938 363134
rect 64022 362898 64258 363134
rect 64342 362898 64578 363134
rect 64662 362898 64898 363134
rect 64982 362898 65218 363134
rect 65302 362898 65538 363134
rect 65622 362898 65858 363134
rect 504050 363218 504286 363454
rect 504370 363218 504606 363454
rect 504690 363218 504926 363454
rect 505010 363218 505246 363454
rect 505330 363218 505566 363454
rect 505650 363218 505886 363454
rect 505970 363218 506206 363454
rect 506290 363218 506526 363454
rect 506610 363218 506846 363454
rect 504050 362898 504286 363134
rect 504370 362898 504606 363134
rect 504690 362898 504926 363134
rect 505010 362898 505246 363134
rect 505330 362898 505566 363134
rect 505650 362898 505886 363134
rect 505970 362898 506206 363134
rect 506290 362898 506526 363134
rect 506610 362898 506846 363134
rect 59062 345218 59298 345454
rect 59382 345218 59618 345454
rect 59702 345218 59938 345454
rect 60022 345218 60258 345454
rect 60342 345218 60578 345454
rect 60662 345218 60898 345454
rect 60982 345218 61218 345454
rect 61302 345218 61538 345454
rect 61622 345218 61858 345454
rect 59062 344898 59298 345134
rect 59382 344898 59618 345134
rect 59702 344898 59938 345134
rect 60022 344898 60258 345134
rect 60342 344898 60578 345134
rect 60662 344898 60898 345134
rect 60982 344898 61218 345134
rect 61302 344898 61538 345134
rect 61622 344898 61858 345134
rect 71177 345218 71413 345454
rect 71177 344898 71413 345134
rect 166241 345218 166477 345454
rect 166241 344898 166477 345134
rect 403133 345218 403369 345454
rect 403133 344898 403369 345134
rect 498197 345218 498433 345454
rect 498197 344898 498433 345134
rect 508050 345218 508286 345454
rect 508370 345218 508606 345454
rect 508690 345218 508926 345454
rect 509010 345218 509246 345454
rect 509330 345218 509566 345454
rect 509650 345218 509886 345454
rect 509970 345218 510206 345454
rect 510290 345218 510526 345454
rect 510610 345218 510846 345454
rect 508050 344898 508286 345134
rect 508370 344898 508606 345134
rect 508690 344898 508926 345134
rect 509010 344898 509246 345134
rect 509330 344898 509566 345134
rect 509650 344898 509886 345134
rect 509970 344898 510206 345134
rect 510290 344898 510526 345134
rect 510610 344898 510846 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 63062 327218 63298 327454
rect 63382 327218 63618 327454
rect 63702 327218 63938 327454
rect 64022 327218 64258 327454
rect 64342 327218 64578 327454
rect 64662 327218 64898 327454
rect 64982 327218 65218 327454
rect 65302 327218 65538 327454
rect 65622 327218 65858 327454
rect 63062 326898 63298 327134
rect 63382 326898 63618 327134
rect 63702 326898 63938 327134
rect 64022 326898 64258 327134
rect 64342 326898 64578 327134
rect 64662 326898 64898 327134
rect 64982 326898 65218 327134
rect 65302 326898 65538 327134
rect 65622 326898 65858 327134
rect 71857 327218 72093 327454
rect 71857 326898 72093 327134
rect 165561 327218 165797 327454
rect 165561 326898 165797 327134
rect 403813 327218 404049 327454
rect 403813 326898 404049 327134
rect 497517 327218 497753 327454
rect 497517 326898 497753 327134
rect 504050 327218 504286 327454
rect 504370 327218 504606 327454
rect 504690 327218 504926 327454
rect 505010 327218 505246 327454
rect 505330 327218 505566 327454
rect 505650 327218 505886 327454
rect 505970 327218 506206 327454
rect 506290 327218 506526 327454
rect 506610 327218 506846 327454
rect 504050 326898 504286 327134
rect 504370 326898 504606 327134
rect 504690 326898 504926 327134
rect 505010 326898 505246 327134
rect 505330 326898 505566 327134
rect 505650 326898 505886 327134
rect 505970 326898 506206 327134
rect 506290 326898 506526 327134
rect 506610 326898 506846 327134
rect 59062 309218 59298 309454
rect 59382 309218 59618 309454
rect 59702 309218 59938 309454
rect 60022 309218 60258 309454
rect 60342 309218 60578 309454
rect 60662 309218 60898 309454
rect 60982 309218 61218 309454
rect 61302 309218 61538 309454
rect 61622 309218 61858 309454
rect 59062 308898 59298 309134
rect 59382 308898 59618 309134
rect 59702 308898 59938 309134
rect 60022 308898 60258 309134
rect 60342 308898 60578 309134
rect 60662 308898 60898 309134
rect 60982 308898 61218 309134
rect 61302 308898 61538 309134
rect 61622 308898 61858 309134
rect 71177 309218 71413 309454
rect 71177 308898 71413 309134
rect 166241 309218 166477 309454
rect 166241 308898 166477 309134
rect 403133 309218 403369 309454
rect 403133 308898 403369 309134
rect 498197 309218 498433 309454
rect 498197 308898 498433 309134
rect 508050 309218 508286 309454
rect 508370 309218 508606 309454
rect 508690 309218 508926 309454
rect 509010 309218 509246 309454
rect 509330 309218 509566 309454
rect 509650 309218 509886 309454
rect 509970 309218 510206 309454
rect 510290 309218 510526 309454
rect 510610 309218 510846 309454
rect 508050 308898 508286 309134
rect 508370 308898 508606 309134
rect 508690 308898 508926 309134
rect 509010 308898 509246 309134
rect 509330 308898 509566 309134
rect 509650 308898 509886 309134
rect 509970 308898 510206 309134
rect 510290 308898 510526 309134
rect 510610 308898 510846 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 63062 291218 63298 291454
rect 63382 291218 63618 291454
rect 63702 291218 63938 291454
rect 64022 291218 64258 291454
rect 64342 291218 64578 291454
rect 64662 291218 64898 291454
rect 64982 291218 65218 291454
rect 65302 291218 65538 291454
rect 65622 291218 65858 291454
rect 63062 290898 63298 291134
rect 63382 290898 63618 291134
rect 63702 290898 63938 291134
rect 64022 290898 64258 291134
rect 64342 290898 64578 291134
rect 64662 290898 64898 291134
rect 64982 290898 65218 291134
rect 65302 290898 65538 291134
rect 65622 290898 65858 291134
rect 71857 291218 72093 291454
rect 71857 290898 72093 291134
rect 165561 291218 165797 291454
rect 165561 290898 165797 291134
rect 403813 291218 404049 291454
rect 403813 290898 404049 291134
rect 497517 291218 497753 291454
rect 497517 290898 497753 291134
rect 504050 291218 504286 291454
rect 504370 291218 504606 291454
rect 504690 291218 504926 291454
rect 505010 291218 505246 291454
rect 505330 291218 505566 291454
rect 505650 291218 505886 291454
rect 505970 291218 506206 291454
rect 506290 291218 506526 291454
rect 506610 291218 506846 291454
rect 504050 290898 504286 291134
rect 504370 290898 504606 291134
rect 504690 290898 504926 291134
rect 505010 290898 505246 291134
rect 505330 290898 505566 291134
rect 505650 290898 505886 291134
rect 505970 290898 506206 291134
rect 506290 290898 506526 291134
rect 506610 290898 506846 291134
rect 59062 273218 59298 273454
rect 59382 273218 59618 273454
rect 59702 273218 59938 273454
rect 60022 273218 60258 273454
rect 60342 273218 60578 273454
rect 60662 273218 60898 273454
rect 60982 273218 61218 273454
rect 61302 273218 61538 273454
rect 61622 273218 61858 273454
rect 59062 272898 59298 273134
rect 59382 272898 59618 273134
rect 59702 272898 59938 273134
rect 60022 272898 60258 273134
rect 60342 272898 60578 273134
rect 60662 272898 60898 273134
rect 60982 272898 61218 273134
rect 61302 272898 61538 273134
rect 61622 272898 61858 273134
rect 508050 273218 508286 273454
rect 508370 273218 508606 273454
rect 508690 273218 508926 273454
rect 509010 273218 509246 273454
rect 509330 273218 509566 273454
rect 509650 273218 509886 273454
rect 509970 273218 510206 273454
rect 510290 273218 510526 273454
rect 510610 273218 510846 273454
rect 508050 272898 508286 273134
rect 508370 272898 508606 273134
rect 508690 272898 508926 273134
rect 509010 272898 509246 273134
rect 509330 272898 509566 273134
rect 509650 272898 509886 273134
rect 509970 272898 510206 273134
rect 510290 272898 510526 273134
rect 510610 272898 510846 273134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 63062 255218 63298 255454
rect 63382 255218 63618 255454
rect 63702 255218 63938 255454
rect 64022 255218 64258 255454
rect 64342 255218 64578 255454
rect 64662 255218 64898 255454
rect 64982 255218 65218 255454
rect 65302 255218 65538 255454
rect 65622 255218 65858 255454
rect 63062 254898 63298 255134
rect 63382 254898 63618 255134
rect 63702 254898 63938 255134
rect 64022 254898 64258 255134
rect 64342 254898 64578 255134
rect 64662 254898 64898 255134
rect 64982 254898 65218 255134
rect 65302 254898 65538 255134
rect 65622 254898 65858 255134
rect 504050 255218 504286 255454
rect 504370 255218 504606 255454
rect 504690 255218 504926 255454
rect 505010 255218 505246 255454
rect 505330 255218 505566 255454
rect 505650 255218 505886 255454
rect 505970 255218 506206 255454
rect 506290 255218 506526 255454
rect 506610 255218 506846 255454
rect 504050 254898 504286 255134
rect 504370 254898 504606 255134
rect 504690 254898 504926 255134
rect 505010 254898 505246 255134
rect 505330 254898 505566 255134
rect 505650 254898 505886 255134
rect 505970 254898 506206 255134
rect 506290 254898 506526 255134
rect 506610 254898 506846 255134
rect 59062 237218 59298 237454
rect 59382 237218 59618 237454
rect 59702 237218 59938 237454
rect 60022 237218 60258 237454
rect 60342 237218 60578 237454
rect 60662 237218 60898 237454
rect 60982 237218 61218 237454
rect 61302 237218 61538 237454
rect 61622 237218 61858 237454
rect 59062 236898 59298 237134
rect 59382 236898 59618 237134
rect 59702 236898 59938 237134
rect 60022 236898 60258 237134
rect 60342 236898 60578 237134
rect 60662 236898 60898 237134
rect 60982 236898 61218 237134
rect 61302 236898 61538 237134
rect 61622 236898 61858 237134
rect 71177 237218 71413 237454
rect 71177 236898 71413 237134
rect 166241 237218 166477 237454
rect 166241 236898 166477 237134
rect 403133 237218 403369 237454
rect 403133 236898 403369 237134
rect 498197 237218 498433 237454
rect 498197 236898 498433 237134
rect 508050 237218 508286 237454
rect 508370 237218 508606 237454
rect 508690 237218 508926 237454
rect 509010 237218 509246 237454
rect 509330 237218 509566 237454
rect 509650 237218 509886 237454
rect 509970 237218 510206 237454
rect 510290 237218 510526 237454
rect 510610 237218 510846 237454
rect 508050 236898 508286 237134
rect 508370 236898 508606 237134
rect 508690 236898 508926 237134
rect 509010 236898 509246 237134
rect 509330 236898 509566 237134
rect 509650 236898 509886 237134
rect 509970 236898 510206 237134
rect 510290 236898 510526 237134
rect 510610 236898 510846 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 63062 219218 63298 219454
rect 63382 219218 63618 219454
rect 63702 219218 63938 219454
rect 64022 219218 64258 219454
rect 64342 219218 64578 219454
rect 64662 219218 64898 219454
rect 64982 219218 65218 219454
rect 65302 219218 65538 219454
rect 65622 219218 65858 219454
rect 63062 218898 63298 219134
rect 63382 218898 63618 219134
rect 63702 218898 63938 219134
rect 64022 218898 64258 219134
rect 64342 218898 64578 219134
rect 64662 218898 64898 219134
rect 64982 218898 65218 219134
rect 65302 218898 65538 219134
rect 65622 218898 65858 219134
rect 71857 219218 72093 219454
rect 71857 218898 72093 219134
rect 165561 219218 165797 219454
rect 165561 218898 165797 219134
rect 403813 219218 404049 219454
rect 403813 218898 404049 219134
rect 497517 219218 497753 219454
rect 497517 218898 497753 219134
rect 504050 219218 504286 219454
rect 504370 219218 504606 219454
rect 504690 219218 504926 219454
rect 505010 219218 505246 219454
rect 505330 219218 505566 219454
rect 505650 219218 505886 219454
rect 505970 219218 506206 219454
rect 506290 219218 506526 219454
rect 506610 219218 506846 219454
rect 504050 218898 504286 219134
rect 504370 218898 504606 219134
rect 504690 218898 504926 219134
rect 505010 218898 505246 219134
rect 505330 218898 505566 219134
rect 505650 218898 505886 219134
rect 505970 218898 506206 219134
rect 506290 218898 506526 219134
rect 506610 218898 506846 219134
rect 59062 201218 59298 201454
rect 59382 201218 59618 201454
rect 59702 201218 59938 201454
rect 60022 201218 60258 201454
rect 60342 201218 60578 201454
rect 60662 201218 60898 201454
rect 60982 201218 61218 201454
rect 61302 201218 61538 201454
rect 61622 201218 61858 201454
rect 59062 200898 59298 201134
rect 59382 200898 59618 201134
rect 59702 200898 59938 201134
rect 60022 200898 60258 201134
rect 60342 200898 60578 201134
rect 60662 200898 60898 201134
rect 60982 200898 61218 201134
rect 61302 200898 61538 201134
rect 61622 200898 61858 201134
rect 71177 201218 71413 201454
rect 71177 200898 71413 201134
rect 166241 201218 166477 201454
rect 166241 200898 166477 201134
rect 403133 201218 403369 201454
rect 403133 200898 403369 201134
rect 498197 201218 498433 201454
rect 498197 200898 498433 201134
rect 508050 201218 508286 201454
rect 508370 201218 508606 201454
rect 508690 201218 508926 201454
rect 509010 201218 509246 201454
rect 509330 201218 509566 201454
rect 509650 201218 509886 201454
rect 509970 201218 510206 201454
rect 510290 201218 510526 201454
rect 510610 201218 510846 201454
rect 508050 200898 508286 201134
rect 508370 200898 508606 201134
rect 508690 200898 508926 201134
rect 509010 200898 509246 201134
rect 509330 200898 509566 201134
rect 509650 200898 509886 201134
rect 509970 200898 510206 201134
rect 510290 200898 510526 201134
rect 510610 200898 510846 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 63062 183218 63298 183454
rect 63382 183218 63618 183454
rect 63702 183218 63938 183454
rect 64022 183218 64258 183454
rect 64342 183218 64578 183454
rect 64662 183218 64898 183454
rect 64982 183218 65218 183454
rect 65302 183218 65538 183454
rect 65622 183218 65858 183454
rect 63062 182898 63298 183134
rect 63382 182898 63618 183134
rect 63702 182898 63938 183134
rect 64022 182898 64258 183134
rect 64342 182898 64578 183134
rect 64662 182898 64898 183134
rect 64982 182898 65218 183134
rect 65302 182898 65538 183134
rect 65622 182898 65858 183134
rect 71857 183218 72093 183454
rect 71857 182898 72093 183134
rect 165561 183218 165797 183454
rect 165561 182898 165797 183134
rect 403813 183218 404049 183454
rect 403813 182898 404049 183134
rect 497517 183218 497753 183454
rect 497517 182898 497753 183134
rect 504050 183218 504286 183454
rect 504370 183218 504606 183454
rect 504690 183218 504926 183454
rect 505010 183218 505246 183454
rect 505330 183218 505566 183454
rect 505650 183218 505886 183454
rect 505970 183218 506206 183454
rect 506290 183218 506526 183454
rect 506610 183218 506846 183454
rect 504050 182898 504286 183134
rect 504370 182898 504606 183134
rect 504690 182898 504926 183134
rect 505010 182898 505246 183134
rect 505330 182898 505566 183134
rect 505650 182898 505886 183134
rect 505970 182898 506206 183134
rect 506290 182898 506526 183134
rect 506610 182898 506846 183134
rect 59062 165218 59298 165454
rect 59382 165218 59618 165454
rect 59702 165218 59938 165454
rect 60022 165218 60258 165454
rect 60342 165218 60578 165454
rect 60662 165218 60898 165454
rect 60982 165218 61218 165454
rect 61302 165218 61538 165454
rect 61622 165218 61858 165454
rect 59062 164898 59298 165134
rect 59382 164898 59618 165134
rect 59702 164898 59938 165134
rect 60022 164898 60258 165134
rect 60342 164898 60578 165134
rect 60662 164898 60898 165134
rect 60982 164898 61218 165134
rect 61302 164898 61538 165134
rect 61622 164898 61858 165134
rect 508050 165218 508286 165454
rect 508370 165218 508606 165454
rect 508690 165218 508926 165454
rect 509010 165218 509246 165454
rect 509330 165218 509566 165454
rect 509650 165218 509886 165454
rect 509970 165218 510206 165454
rect 510290 165218 510526 165454
rect 510610 165218 510846 165454
rect 508050 164898 508286 165134
rect 508370 164898 508606 165134
rect 508690 164898 508926 165134
rect 509010 164898 509246 165134
rect 509330 164898 509566 165134
rect 509650 164898 509886 165134
rect 509970 164898 510206 165134
rect 510290 164898 510526 165134
rect 510610 164898 510846 165134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 63062 147218 63298 147454
rect 63382 147218 63618 147454
rect 63702 147218 63938 147454
rect 64022 147218 64258 147454
rect 64342 147218 64578 147454
rect 64662 147218 64898 147454
rect 64982 147218 65218 147454
rect 65302 147218 65538 147454
rect 65622 147218 65858 147454
rect 63062 146898 63298 147134
rect 63382 146898 63618 147134
rect 63702 146898 63938 147134
rect 64022 146898 64258 147134
rect 64342 146898 64578 147134
rect 64662 146898 64898 147134
rect 64982 146898 65218 147134
rect 65302 146898 65538 147134
rect 65622 146898 65858 147134
rect 71857 147218 72093 147454
rect 71857 146898 72093 147134
rect 165561 147218 165797 147454
rect 165561 146898 165797 147134
rect 403813 147218 404049 147454
rect 403813 146898 404049 147134
rect 497517 147218 497753 147454
rect 497517 146898 497753 147134
rect 504050 147218 504286 147454
rect 504370 147218 504606 147454
rect 504690 147218 504926 147454
rect 505010 147218 505246 147454
rect 505330 147218 505566 147454
rect 505650 147218 505886 147454
rect 505970 147218 506206 147454
rect 506290 147218 506526 147454
rect 506610 147218 506846 147454
rect 504050 146898 504286 147134
rect 504370 146898 504606 147134
rect 504690 146898 504926 147134
rect 505010 146898 505246 147134
rect 505330 146898 505566 147134
rect 505650 146898 505886 147134
rect 505970 146898 506206 147134
rect 506290 146898 506526 147134
rect 506610 146898 506846 147134
rect 59062 129218 59298 129454
rect 59382 129218 59618 129454
rect 59702 129218 59938 129454
rect 60022 129218 60258 129454
rect 60342 129218 60578 129454
rect 60662 129218 60898 129454
rect 60982 129218 61218 129454
rect 61302 129218 61538 129454
rect 61622 129218 61858 129454
rect 59062 128898 59298 129134
rect 59382 128898 59618 129134
rect 59702 128898 59938 129134
rect 60022 128898 60258 129134
rect 60342 128898 60578 129134
rect 60662 128898 60898 129134
rect 60982 128898 61218 129134
rect 61302 128898 61538 129134
rect 61622 128898 61858 129134
rect 71177 129218 71413 129454
rect 71177 128898 71413 129134
rect 166241 129218 166477 129454
rect 166241 128898 166477 129134
rect 403133 129218 403369 129454
rect 403133 128898 403369 129134
rect 498197 129218 498433 129454
rect 498197 128898 498433 129134
rect 508050 129218 508286 129454
rect 508370 129218 508606 129454
rect 508690 129218 508926 129454
rect 509010 129218 509246 129454
rect 509330 129218 509566 129454
rect 509650 129218 509886 129454
rect 509970 129218 510206 129454
rect 510290 129218 510526 129454
rect 510610 129218 510846 129454
rect 508050 128898 508286 129134
rect 508370 128898 508606 129134
rect 508690 128898 508926 129134
rect 509010 128898 509246 129134
rect 509330 128898 509566 129134
rect 509650 128898 509886 129134
rect 509970 128898 510206 129134
rect 510290 128898 510526 129134
rect 510610 128898 510846 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 63062 111218 63298 111454
rect 63382 111218 63618 111454
rect 63702 111218 63938 111454
rect 64022 111218 64258 111454
rect 64342 111218 64578 111454
rect 64662 111218 64898 111454
rect 64982 111218 65218 111454
rect 65302 111218 65538 111454
rect 65622 111218 65858 111454
rect 63062 110898 63298 111134
rect 63382 110898 63618 111134
rect 63702 110898 63938 111134
rect 64022 110898 64258 111134
rect 64342 110898 64578 111134
rect 64662 110898 64898 111134
rect 64982 110898 65218 111134
rect 65302 110898 65538 111134
rect 65622 110898 65858 111134
rect 71857 111218 72093 111454
rect 71857 110898 72093 111134
rect 165561 111218 165797 111454
rect 165561 110898 165797 111134
rect 403813 111218 404049 111454
rect 403813 110898 404049 111134
rect 497517 111218 497753 111454
rect 497517 110898 497753 111134
rect 504050 111218 504286 111454
rect 504370 111218 504606 111454
rect 504690 111218 504926 111454
rect 505010 111218 505246 111454
rect 505330 111218 505566 111454
rect 505650 111218 505886 111454
rect 505970 111218 506206 111454
rect 506290 111218 506526 111454
rect 506610 111218 506846 111454
rect 504050 110898 504286 111134
rect 504370 110898 504606 111134
rect 504690 110898 504926 111134
rect 505010 110898 505246 111134
rect 505330 110898 505566 111134
rect 505650 110898 505886 111134
rect 505970 110898 506206 111134
rect 506290 110898 506526 111134
rect 506610 110898 506846 111134
rect 59062 93218 59298 93454
rect 59382 93218 59618 93454
rect 59702 93218 59938 93454
rect 60022 93218 60258 93454
rect 60342 93218 60578 93454
rect 60662 93218 60898 93454
rect 60982 93218 61218 93454
rect 61302 93218 61538 93454
rect 61622 93218 61858 93454
rect 59062 92898 59298 93134
rect 59382 92898 59618 93134
rect 59702 92898 59938 93134
rect 60022 92898 60258 93134
rect 60342 92898 60578 93134
rect 60662 92898 60898 93134
rect 60982 92898 61218 93134
rect 61302 92898 61538 93134
rect 61622 92898 61858 93134
rect 71177 93218 71413 93454
rect 71177 92898 71413 93134
rect 166241 93218 166477 93454
rect 166241 92898 166477 93134
rect 403133 93218 403369 93454
rect 403133 92898 403369 93134
rect 498197 93218 498433 93454
rect 498197 92898 498433 93134
rect 508050 93218 508286 93454
rect 508370 93218 508606 93454
rect 508690 93218 508926 93454
rect 509010 93218 509246 93454
rect 509330 93218 509566 93454
rect 509650 93218 509886 93454
rect 509970 93218 510206 93454
rect 510290 93218 510526 93454
rect 510610 93218 510846 93454
rect 508050 92898 508286 93134
rect 508370 92898 508606 93134
rect 508690 92898 508926 93134
rect 509010 92898 509246 93134
rect 509330 92898 509566 93134
rect 509650 92898 509886 93134
rect 509970 92898 510206 93134
rect 510290 92898 510526 93134
rect 510610 92898 510846 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 63062 75218 63298 75454
rect 63382 75218 63618 75454
rect 63702 75218 63938 75454
rect 64022 75218 64258 75454
rect 64342 75218 64578 75454
rect 64662 75218 64898 75454
rect 64982 75218 65218 75454
rect 65302 75218 65538 75454
rect 65622 75218 65858 75454
rect 63062 74898 63298 75134
rect 63382 74898 63618 75134
rect 63702 74898 63938 75134
rect 64022 74898 64258 75134
rect 64342 74898 64578 75134
rect 64662 74898 64898 75134
rect 64982 74898 65218 75134
rect 65302 74898 65538 75134
rect 65622 74898 65858 75134
rect 504050 75218 504286 75454
rect 504370 75218 504606 75454
rect 504690 75218 504926 75454
rect 505010 75218 505246 75454
rect 505330 75218 505566 75454
rect 505650 75218 505886 75454
rect 505970 75218 506206 75454
rect 506290 75218 506526 75454
rect 506610 75218 506846 75454
rect 504050 74898 504286 75134
rect 504370 74898 504606 75134
rect 504690 74898 504926 75134
rect 505010 74898 505246 75134
rect 505330 74898 505566 75134
rect 505650 74898 505886 75134
rect 505970 74898 506206 75134
rect 506290 74898 506526 75134
rect 506610 74898 506846 75134
rect 59062 57218 59298 57454
rect 59382 57218 59618 57454
rect 59702 57218 59938 57454
rect 60022 57218 60258 57454
rect 60342 57218 60578 57454
rect 60662 57218 60898 57454
rect 60982 57218 61218 57454
rect 61302 57218 61538 57454
rect 61622 57218 61858 57454
rect 59062 56898 59298 57134
rect 59382 56898 59618 57134
rect 59702 56898 59938 57134
rect 60022 56898 60258 57134
rect 60342 56898 60578 57134
rect 60662 56898 60898 57134
rect 60982 56898 61218 57134
rect 61302 56898 61538 57134
rect 61622 56898 61858 57134
rect 508050 57218 508286 57454
rect 508370 57218 508606 57454
rect 508690 57218 508926 57454
rect 509010 57218 509246 57454
rect 509330 57218 509566 57454
rect 509650 57218 509886 57454
rect 509970 57218 510206 57454
rect 510290 57218 510526 57454
rect 510610 57218 510846 57454
rect 508050 56898 508286 57134
rect 508370 56898 508606 57134
rect 508690 56898 508926 57134
rect 509010 56898 509246 57134
rect 509330 56898 509566 57134
rect 509650 56898 509886 57134
rect 509970 56898 510206 57134
rect 510290 56898 510526 57134
rect 510610 56898 510846 57134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 63062 39218 63298 39454
rect 63382 39218 63618 39454
rect 63702 39218 63938 39454
rect 64022 39218 64258 39454
rect 64342 39218 64578 39454
rect 64662 39218 64898 39454
rect 64982 39218 65218 39454
rect 65302 39218 65538 39454
rect 65622 39218 65858 39454
rect 63062 38898 63298 39134
rect 63382 38898 63618 39134
rect 63702 38898 63938 39134
rect 64022 38898 64258 39134
rect 64342 38898 64578 39134
rect 64662 38898 64898 39134
rect 64982 38898 65218 39134
rect 65302 38898 65538 39134
rect 65622 38898 65858 39134
rect 504050 39218 504286 39454
rect 504370 39218 504606 39454
rect 504690 39218 504926 39454
rect 505010 39218 505246 39454
rect 505330 39218 505566 39454
rect 505650 39218 505886 39454
rect 505970 39218 506206 39454
rect 506290 39218 506526 39454
rect 506610 39218 506846 39454
rect 504050 38898 504286 39134
rect 504370 38898 504606 39134
rect 504690 38898 504926 39134
rect 505010 38898 505246 39134
rect 505330 38898 505566 39134
rect 505650 38898 505886 39134
rect 505970 38898 506206 39134
rect 506290 38898 506526 39134
rect 506610 38898 506846 39134
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 59062 453454
rect 59298 453218 59382 453454
rect 59618 453218 59702 453454
rect 59938 453218 60022 453454
rect 60258 453218 60342 453454
rect 60578 453218 60662 453454
rect 60898 453218 60982 453454
rect 61218 453218 61302 453454
rect 61538 453218 61622 453454
rect 61858 453218 71177 453454
rect 71413 453218 166241 453454
rect 166477 453218 403133 453454
rect 403369 453218 498197 453454
rect 498433 453218 508050 453454
rect 508286 453218 508370 453454
rect 508606 453218 508690 453454
rect 508926 453218 509010 453454
rect 509246 453218 509330 453454
rect 509566 453218 509650 453454
rect 509886 453218 509970 453454
rect 510206 453218 510290 453454
rect 510526 453218 510610 453454
rect 510846 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 59062 453134
rect 59298 452898 59382 453134
rect 59618 452898 59702 453134
rect 59938 452898 60022 453134
rect 60258 452898 60342 453134
rect 60578 452898 60662 453134
rect 60898 452898 60982 453134
rect 61218 452898 61302 453134
rect 61538 452898 61622 453134
rect 61858 452898 71177 453134
rect 71413 452898 166241 453134
rect 166477 452898 403133 453134
rect 403369 452898 498197 453134
rect 498433 452898 508050 453134
rect 508286 452898 508370 453134
rect 508606 452898 508690 453134
rect 508926 452898 509010 453134
rect 509246 452898 509330 453134
rect 509566 452898 509650 453134
rect 509886 452898 509970 453134
rect 510206 452898 510290 453134
rect 510526 452898 510610 453134
rect 510846 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 63062 435454
rect 63298 435218 63382 435454
rect 63618 435218 63702 435454
rect 63938 435218 64022 435454
rect 64258 435218 64342 435454
rect 64578 435218 64662 435454
rect 64898 435218 64982 435454
rect 65218 435218 65302 435454
rect 65538 435218 65622 435454
rect 65858 435218 71857 435454
rect 72093 435218 165561 435454
rect 165797 435218 403813 435454
rect 404049 435218 497517 435454
rect 497753 435218 504050 435454
rect 504286 435218 504370 435454
rect 504606 435218 504690 435454
rect 504926 435218 505010 435454
rect 505246 435218 505330 435454
rect 505566 435218 505650 435454
rect 505886 435218 505970 435454
rect 506206 435218 506290 435454
rect 506526 435218 506610 435454
rect 506846 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 63062 435134
rect 63298 434898 63382 435134
rect 63618 434898 63702 435134
rect 63938 434898 64022 435134
rect 64258 434898 64342 435134
rect 64578 434898 64662 435134
rect 64898 434898 64982 435134
rect 65218 434898 65302 435134
rect 65538 434898 65622 435134
rect 65858 434898 71857 435134
rect 72093 434898 165561 435134
rect 165797 434898 403813 435134
rect 404049 434898 497517 435134
rect 497753 434898 504050 435134
rect 504286 434898 504370 435134
rect 504606 434898 504690 435134
rect 504926 434898 505010 435134
rect 505246 434898 505330 435134
rect 505566 434898 505650 435134
rect 505886 434898 505970 435134
rect 506206 434898 506290 435134
rect 506526 434898 506610 435134
rect 506846 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 59062 417454
rect 59298 417218 59382 417454
rect 59618 417218 59702 417454
rect 59938 417218 60022 417454
rect 60258 417218 60342 417454
rect 60578 417218 60662 417454
rect 60898 417218 60982 417454
rect 61218 417218 61302 417454
rect 61538 417218 61622 417454
rect 61858 417218 71177 417454
rect 71413 417218 166241 417454
rect 166477 417218 403133 417454
rect 403369 417218 498197 417454
rect 498433 417218 508050 417454
rect 508286 417218 508370 417454
rect 508606 417218 508690 417454
rect 508926 417218 509010 417454
rect 509246 417218 509330 417454
rect 509566 417218 509650 417454
rect 509886 417218 509970 417454
rect 510206 417218 510290 417454
rect 510526 417218 510610 417454
rect 510846 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 59062 417134
rect 59298 416898 59382 417134
rect 59618 416898 59702 417134
rect 59938 416898 60022 417134
rect 60258 416898 60342 417134
rect 60578 416898 60662 417134
rect 60898 416898 60982 417134
rect 61218 416898 61302 417134
rect 61538 416898 61622 417134
rect 61858 416898 71177 417134
rect 71413 416898 166241 417134
rect 166477 416898 403133 417134
rect 403369 416898 498197 417134
rect 498433 416898 508050 417134
rect 508286 416898 508370 417134
rect 508606 416898 508690 417134
rect 508926 416898 509010 417134
rect 509246 416898 509330 417134
rect 509566 416898 509650 417134
rect 509886 416898 509970 417134
rect 510206 416898 510290 417134
rect 510526 416898 510610 417134
rect 510846 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 63062 399454
rect 63298 399218 63382 399454
rect 63618 399218 63702 399454
rect 63938 399218 64022 399454
rect 64258 399218 64342 399454
rect 64578 399218 64662 399454
rect 64898 399218 64982 399454
rect 65218 399218 65302 399454
rect 65538 399218 65622 399454
rect 65858 399218 71857 399454
rect 72093 399218 165561 399454
rect 165797 399218 403813 399454
rect 404049 399218 497517 399454
rect 497753 399218 504050 399454
rect 504286 399218 504370 399454
rect 504606 399218 504690 399454
rect 504926 399218 505010 399454
rect 505246 399218 505330 399454
rect 505566 399218 505650 399454
rect 505886 399218 505970 399454
rect 506206 399218 506290 399454
rect 506526 399218 506610 399454
rect 506846 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 63062 399134
rect 63298 398898 63382 399134
rect 63618 398898 63702 399134
rect 63938 398898 64022 399134
rect 64258 398898 64342 399134
rect 64578 398898 64662 399134
rect 64898 398898 64982 399134
rect 65218 398898 65302 399134
rect 65538 398898 65622 399134
rect 65858 398898 71857 399134
rect 72093 398898 165561 399134
rect 165797 398898 403813 399134
rect 404049 398898 497517 399134
rect 497753 398898 504050 399134
rect 504286 398898 504370 399134
rect 504606 398898 504690 399134
rect 504926 398898 505010 399134
rect 505246 398898 505330 399134
rect 505566 398898 505650 399134
rect 505886 398898 505970 399134
rect 506206 398898 506290 399134
rect 506526 398898 506610 399134
rect 506846 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 59062 381454
rect 59298 381218 59382 381454
rect 59618 381218 59702 381454
rect 59938 381218 60022 381454
rect 60258 381218 60342 381454
rect 60578 381218 60662 381454
rect 60898 381218 60982 381454
rect 61218 381218 61302 381454
rect 61538 381218 61622 381454
rect 61858 381218 71177 381454
rect 71413 381218 166241 381454
rect 166477 381218 403133 381454
rect 403369 381218 498197 381454
rect 498433 381218 508050 381454
rect 508286 381218 508370 381454
rect 508606 381218 508690 381454
rect 508926 381218 509010 381454
rect 509246 381218 509330 381454
rect 509566 381218 509650 381454
rect 509886 381218 509970 381454
rect 510206 381218 510290 381454
rect 510526 381218 510610 381454
rect 510846 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 59062 381134
rect 59298 380898 59382 381134
rect 59618 380898 59702 381134
rect 59938 380898 60022 381134
rect 60258 380898 60342 381134
rect 60578 380898 60662 381134
rect 60898 380898 60982 381134
rect 61218 380898 61302 381134
rect 61538 380898 61622 381134
rect 61858 380898 71177 381134
rect 71413 380898 166241 381134
rect 166477 380898 403133 381134
rect 403369 380898 498197 381134
rect 498433 380898 508050 381134
rect 508286 380898 508370 381134
rect 508606 380898 508690 381134
rect 508926 380898 509010 381134
rect 509246 380898 509330 381134
rect 509566 380898 509650 381134
rect 509886 380898 509970 381134
rect 510206 380898 510290 381134
rect 510526 380898 510610 381134
rect 510846 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 63062 363454
rect 63298 363218 63382 363454
rect 63618 363218 63702 363454
rect 63938 363218 64022 363454
rect 64258 363218 64342 363454
rect 64578 363218 64662 363454
rect 64898 363218 64982 363454
rect 65218 363218 65302 363454
rect 65538 363218 65622 363454
rect 65858 363218 504050 363454
rect 504286 363218 504370 363454
rect 504606 363218 504690 363454
rect 504926 363218 505010 363454
rect 505246 363218 505330 363454
rect 505566 363218 505650 363454
rect 505886 363218 505970 363454
rect 506206 363218 506290 363454
rect 506526 363218 506610 363454
rect 506846 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 63062 363134
rect 63298 362898 63382 363134
rect 63618 362898 63702 363134
rect 63938 362898 64022 363134
rect 64258 362898 64342 363134
rect 64578 362898 64662 363134
rect 64898 362898 64982 363134
rect 65218 362898 65302 363134
rect 65538 362898 65622 363134
rect 65858 362898 504050 363134
rect 504286 362898 504370 363134
rect 504606 362898 504690 363134
rect 504926 362898 505010 363134
rect 505246 362898 505330 363134
rect 505566 362898 505650 363134
rect 505886 362898 505970 363134
rect 506206 362898 506290 363134
rect 506526 362898 506610 363134
rect 506846 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 59062 345454
rect 59298 345218 59382 345454
rect 59618 345218 59702 345454
rect 59938 345218 60022 345454
rect 60258 345218 60342 345454
rect 60578 345218 60662 345454
rect 60898 345218 60982 345454
rect 61218 345218 61302 345454
rect 61538 345218 61622 345454
rect 61858 345218 71177 345454
rect 71413 345218 166241 345454
rect 166477 345218 403133 345454
rect 403369 345218 498197 345454
rect 498433 345218 508050 345454
rect 508286 345218 508370 345454
rect 508606 345218 508690 345454
rect 508926 345218 509010 345454
rect 509246 345218 509330 345454
rect 509566 345218 509650 345454
rect 509886 345218 509970 345454
rect 510206 345218 510290 345454
rect 510526 345218 510610 345454
rect 510846 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 59062 345134
rect 59298 344898 59382 345134
rect 59618 344898 59702 345134
rect 59938 344898 60022 345134
rect 60258 344898 60342 345134
rect 60578 344898 60662 345134
rect 60898 344898 60982 345134
rect 61218 344898 61302 345134
rect 61538 344898 61622 345134
rect 61858 344898 71177 345134
rect 71413 344898 166241 345134
rect 166477 344898 403133 345134
rect 403369 344898 498197 345134
rect 498433 344898 508050 345134
rect 508286 344898 508370 345134
rect 508606 344898 508690 345134
rect 508926 344898 509010 345134
rect 509246 344898 509330 345134
rect 509566 344898 509650 345134
rect 509886 344898 509970 345134
rect 510206 344898 510290 345134
rect 510526 344898 510610 345134
rect 510846 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 63062 327454
rect 63298 327218 63382 327454
rect 63618 327218 63702 327454
rect 63938 327218 64022 327454
rect 64258 327218 64342 327454
rect 64578 327218 64662 327454
rect 64898 327218 64982 327454
rect 65218 327218 65302 327454
rect 65538 327218 65622 327454
rect 65858 327218 71857 327454
rect 72093 327218 165561 327454
rect 165797 327218 403813 327454
rect 404049 327218 497517 327454
rect 497753 327218 504050 327454
rect 504286 327218 504370 327454
rect 504606 327218 504690 327454
rect 504926 327218 505010 327454
rect 505246 327218 505330 327454
rect 505566 327218 505650 327454
rect 505886 327218 505970 327454
rect 506206 327218 506290 327454
rect 506526 327218 506610 327454
rect 506846 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 63062 327134
rect 63298 326898 63382 327134
rect 63618 326898 63702 327134
rect 63938 326898 64022 327134
rect 64258 326898 64342 327134
rect 64578 326898 64662 327134
rect 64898 326898 64982 327134
rect 65218 326898 65302 327134
rect 65538 326898 65622 327134
rect 65858 326898 71857 327134
rect 72093 326898 165561 327134
rect 165797 326898 403813 327134
rect 404049 326898 497517 327134
rect 497753 326898 504050 327134
rect 504286 326898 504370 327134
rect 504606 326898 504690 327134
rect 504926 326898 505010 327134
rect 505246 326898 505330 327134
rect 505566 326898 505650 327134
rect 505886 326898 505970 327134
rect 506206 326898 506290 327134
rect 506526 326898 506610 327134
rect 506846 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 59062 309454
rect 59298 309218 59382 309454
rect 59618 309218 59702 309454
rect 59938 309218 60022 309454
rect 60258 309218 60342 309454
rect 60578 309218 60662 309454
rect 60898 309218 60982 309454
rect 61218 309218 61302 309454
rect 61538 309218 61622 309454
rect 61858 309218 71177 309454
rect 71413 309218 166241 309454
rect 166477 309218 403133 309454
rect 403369 309218 498197 309454
rect 498433 309218 508050 309454
rect 508286 309218 508370 309454
rect 508606 309218 508690 309454
rect 508926 309218 509010 309454
rect 509246 309218 509330 309454
rect 509566 309218 509650 309454
rect 509886 309218 509970 309454
rect 510206 309218 510290 309454
rect 510526 309218 510610 309454
rect 510846 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 59062 309134
rect 59298 308898 59382 309134
rect 59618 308898 59702 309134
rect 59938 308898 60022 309134
rect 60258 308898 60342 309134
rect 60578 308898 60662 309134
rect 60898 308898 60982 309134
rect 61218 308898 61302 309134
rect 61538 308898 61622 309134
rect 61858 308898 71177 309134
rect 71413 308898 166241 309134
rect 166477 308898 403133 309134
rect 403369 308898 498197 309134
rect 498433 308898 508050 309134
rect 508286 308898 508370 309134
rect 508606 308898 508690 309134
rect 508926 308898 509010 309134
rect 509246 308898 509330 309134
rect 509566 308898 509650 309134
rect 509886 308898 509970 309134
rect 510206 308898 510290 309134
rect 510526 308898 510610 309134
rect 510846 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 63062 291454
rect 63298 291218 63382 291454
rect 63618 291218 63702 291454
rect 63938 291218 64022 291454
rect 64258 291218 64342 291454
rect 64578 291218 64662 291454
rect 64898 291218 64982 291454
rect 65218 291218 65302 291454
rect 65538 291218 65622 291454
rect 65858 291218 71857 291454
rect 72093 291218 165561 291454
rect 165797 291218 403813 291454
rect 404049 291218 497517 291454
rect 497753 291218 504050 291454
rect 504286 291218 504370 291454
rect 504606 291218 504690 291454
rect 504926 291218 505010 291454
rect 505246 291218 505330 291454
rect 505566 291218 505650 291454
rect 505886 291218 505970 291454
rect 506206 291218 506290 291454
rect 506526 291218 506610 291454
rect 506846 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 63062 291134
rect 63298 290898 63382 291134
rect 63618 290898 63702 291134
rect 63938 290898 64022 291134
rect 64258 290898 64342 291134
rect 64578 290898 64662 291134
rect 64898 290898 64982 291134
rect 65218 290898 65302 291134
rect 65538 290898 65622 291134
rect 65858 290898 71857 291134
rect 72093 290898 165561 291134
rect 165797 290898 403813 291134
rect 404049 290898 497517 291134
rect 497753 290898 504050 291134
rect 504286 290898 504370 291134
rect 504606 290898 504690 291134
rect 504926 290898 505010 291134
rect 505246 290898 505330 291134
rect 505566 290898 505650 291134
rect 505886 290898 505970 291134
rect 506206 290898 506290 291134
rect 506526 290898 506610 291134
rect 506846 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 59062 273454
rect 59298 273218 59382 273454
rect 59618 273218 59702 273454
rect 59938 273218 60022 273454
rect 60258 273218 60342 273454
rect 60578 273218 60662 273454
rect 60898 273218 60982 273454
rect 61218 273218 61302 273454
rect 61538 273218 61622 273454
rect 61858 273218 508050 273454
rect 508286 273218 508370 273454
rect 508606 273218 508690 273454
rect 508926 273218 509010 273454
rect 509246 273218 509330 273454
rect 509566 273218 509650 273454
rect 509886 273218 509970 273454
rect 510206 273218 510290 273454
rect 510526 273218 510610 273454
rect 510846 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 59062 273134
rect 59298 272898 59382 273134
rect 59618 272898 59702 273134
rect 59938 272898 60022 273134
rect 60258 272898 60342 273134
rect 60578 272898 60662 273134
rect 60898 272898 60982 273134
rect 61218 272898 61302 273134
rect 61538 272898 61622 273134
rect 61858 272898 508050 273134
rect 508286 272898 508370 273134
rect 508606 272898 508690 273134
rect 508926 272898 509010 273134
rect 509246 272898 509330 273134
rect 509566 272898 509650 273134
rect 509886 272898 509970 273134
rect 510206 272898 510290 273134
rect 510526 272898 510610 273134
rect 510846 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 63062 255454
rect 63298 255218 63382 255454
rect 63618 255218 63702 255454
rect 63938 255218 64022 255454
rect 64258 255218 64342 255454
rect 64578 255218 64662 255454
rect 64898 255218 64982 255454
rect 65218 255218 65302 255454
rect 65538 255218 65622 255454
rect 65858 255218 504050 255454
rect 504286 255218 504370 255454
rect 504606 255218 504690 255454
rect 504926 255218 505010 255454
rect 505246 255218 505330 255454
rect 505566 255218 505650 255454
rect 505886 255218 505970 255454
rect 506206 255218 506290 255454
rect 506526 255218 506610 255454
rect 506846 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 63062 255134
rect 63298 254898 63382 255134
rect 63618 254898 63702 255134
rect 63938 254898 64022 255134
rect 64258 254898 64342 255134
rect 64578 254898 64662 255134
rect 64898 254898 64982 255134
rect 65218 254898 65302 255134
rect 65538 254898 65622 255134
rect 65858 254898 504050 255134
rect 504286 254898 504370 255134
rect 504606 254898 504690 255134
rect 504926 254898 505010 255134
rect 505246 254898 505330 255134
rect 505566 254898 505650 255134
rect 505886 254898 505970 255134
rect 506206 254898 506290 255134
rect 506526 254898 506610 255134
rect 506846 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 59062 237454
rect 59298 237218 59382 237454
rect 59618 237218 59702 237454
rect 59938 237218 60022 237454
rect 60258 237218 60342 237454
rect 60578 237218 60662 237454
rect 60898 237218 60982 237454
rect 61218 237218 61302 237454
rect 61538 237218 61622 237454
rect 61858 237218 71177 237454
rect 71413 237218 166241 237454
rect 166477 237218 403133 237454
rect 403369 237218 498197 237454
rect 498433 237218 508050 237454
rect 508286 237218 508370 237454
rect 508606 237218 508690 237454
rect 508926 237218 509010 237454
rect 509246 237218 509330 237454
rect 509566 237218 509650 237454
rect 509886 237218 509970 237454
rect 510206 237218 510290 237454
rect 510526 237218 510610 237454
rect 510846 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 59062 237134
rect 59298 236898 59382 237134
rect 59618 236898 59702 237134
rect 59938 236898 60022 237134
rect 60258 236898 60342 237134
rect 60578 236898 60662 237134
rect 60898 236898 60982 237134
rect 61218 236898 61302 237134
rect 61538 236898 61622 237134
rect 61858 236898 71177 237134
rect 71413 236898 166241 237134
rect 166477 236898 403133 237134
rect 403369 236898 498197 237134
rect 498433 236898 508050 237134
rect 508286 236898 508370 237134
rect 508606 236898 508690 237134
rect 508926 236898 509010 237134
rect 509246 236898 509330 237134
rect 509566 236898 509650 237134
rect 509886 236898 509970 237134
rect 510206 236898 510290 237134
rect 510526 236898 510610 237134
rect 510846 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 63062 219454
rect 63298 219218 63382 219454
rect 63618 219218 63702 219454
rect 63938 219218 64022 219454
rect 64258 219218 64342 219454
rect 64578 219218 64662 219454
rect 64898 219218 64982 219454
rect 65218 219218 65302 219454
rect 65538 219218 65622 219454
rect 65858 219218 71857 219454
rect 72093 219218 165561 219454
rect 165797 219218 403813 219454
rect 404049 219218 497517 219454
rect 497753 219218 504050 219454
rect 504286 219218 504370 219454
rect 504606 219218 504690 219454
rect 504926 219218 505010 219454
rect 505246 219218 505330 219454
rect 505566 219218 505650 219454
rect 505886 219218 505970 219454
rect 506206 219218 506290 219454
rect 506526 219218 506610 219454
rect 506846 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 63062 219134
rect 63298 218898 63382 219134
rect 63618 218898 63702 219134
rect 63938 218898 64022 219134
rect 64258 218898 64342 219134
rect 64578 218898 64662 219134
rect 64898 218898 64982 219134
rect 65218 218898 65302 219134
rect 65538 218898 65622 219134
rect 65858 218898 71857 219134
rect 72093 218898 165561 219134
rect 165797 218898 403813 219134
rect 404049 218898 497517 219134
rect 497753 218898 504050 219134
rect 504286 218898 504370 219134
rect 504606 218898 504690 219134
rect 504926 218898 505010 219134
rect 505246 218898 505330 219134
rect 505566 218898 505650 219134
rect 505886 218898 505970 219134
rect 506206 218898 506290 219134
rect 506526 218898 506610 219134
rect 506846 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 59062 201454
rect 59298 201218 59382 201454
rect 59618 201218 59702 201454
rect 59938 201218 60022 201454
rect 60258 201218 60342 201454
rect 60578 201218 60662 201454
rect 60898 201218 60982 201454
rect 61218 201218 61302 201454
rect 61538 201218 61622 201454
rect 61858 201218 71177 201454
rect 71413 201218 166241 201454
rect 166477 201218 403133 201454
rect 403369 201218 498197 201454
rect 498433 201218 508050 201454
rect 508286 201218 508370 201454
rect 508606 201218 508690 201454
rect 508926 201218 509010 201454
rect 509246 201218 509330 201454
rect 509566 201218 509650 201454
rect 509886 201218 509970 201454
rect 510206 201218 510290 201454
rect 510526 201218 510610 201454
rect 510846 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 59062 201134
rect 59298 200898 59382 201134
rect 59618 200898 59702 201134
rect 59938 200898 60022 201134
rect 60258 200898 60342 201134
rect 60578 200898 60662 201134
rect 60898 200898 60982 201134
rect 61218 200898 61302 201134
rect 61538 200898 61622 201134
rect 61858 200898 71177 201134
rect 71413 200898 166241 201134
rect 166477 200898 403133 201134
rect 403369 200898 498197 201134
rect 498433 200898 508050 201134
rect 508286 200898 508370 201134
rect 508606 200898 508690 201134
rect 508926 200898 509010 201134
rect 509246 200898 509330 201134
rect 509566 200898 509650 201134
rect 509886 200898 509970 201134
rect 510206 200898 510290 201134
rect 510526 200898 510610 201134
rect 510846 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 63062 183454
rect 63298 183218 63382 183454
rect 63618 183218 63702 183454
rect 63938 183218 64022 183454
rect 64258 183218 64342 183454
rect 64578 183218 64662 183454
rect 64898 183218 64982 183454
rect 65218 183218 65302 183454
rect 65538 183218 65622 183454
rect 65858 183218 71857 183454
rect 72093 183218 165561 183454
rect 165797 183218 403813 183454
rect 404049 183218 497517 183454
rect 497753 183218 504050 183454
rect 504286 183218 504370 183454
rect 504606 183218 504690 183454
rect 504926 183218 505010 183454
rect 505246 183218 505330 183454
rect 505566 183218 505650 183454
rect 505886 183218 505970 183454
rect 506206 183218 506290 183454
rect 506526 183218 506610 183454
rect 506846 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 63062 183134
rect 63298 182898 63382 183134
rect 63618 182898 63702 183134
rect 63938 182898 64022 183134
rect 64258 182898 64342 183134
rect 64578 182898 64662 183134
rect 64898 182898 64982 183134
rect 65218 182898 65302 183134
rect 65538 182898 65622 183134
rect 65858 182898 71857 183134
rect 72093 182898 165561 183134
rect 165797 182898 403813 183134
rect 404049 182898 497517 183134
rect 497753 182898 504050 183134
rect 504286 182898 504370 183134
rect 504606 182898 504690 183134
rect 504926 182898 505010 183134
rect 505246 182898 505330 183134
rect 505566 182898 505650 183134
rect 505886 182898 505970 183134
rect 506206 182898 506290 183134
rect 506526 182898 506610 183134
rect 506846 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 59062 165454
rect 59298 165218 59382 165454
rect 59618 165218 59702 165454
rect 59938 165218 60022 165454
rect 60258 165218 60342 165454
rect 60578 165218 60662 165454
rect 60898 165218 60982 165454
rect 61218 165218 61302 165454
rect 61538 165218 61622 165454
rect 61858 165218 508050 165454
rect 508286 165218 508370 165454
rect 508606 165218 508690 165454
rect 508926 165218 509010 165454
rect 509246 165218 509330 165454
rect 509566 165218 509650 165454
rect 509886 165218 509970 165454
rect 510206 165218 510290 165454
rect 510526 165218 510610 165454
rect 510846 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 59062 165134
rect 59298 164898 59382 165134
rect 59618 164898 59702 165134
rect 59938 164898 60022 165134
rect 60258 164898 60342 165134
rect 60578 164898 60662 165134
rect 60898 164898 60982 165134
rect 61218 164898 61302 165134
rect 61538 164898 61622 165134
rect 61858 164898 508050 165134
rect 508286 164898 508370 165134
rect 508606 164898 508690 165134
rect 508926 164898 509010 165134
rect 509246 164898 509330 165134
rect 509566 164898 509650 165134
rect 509886 164898 509970 165134
rect 510206 164898 510290 165134
rect 510526 164898 510610 165134
rect 510846 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 63062 147454
rect 63298 147218 63382 147454
rect 63618 147218 63702 147454
rect 63938 147218 64022 147454
rect 64258 147218 64342 147454
rect 64578 147218 64662 147454
rect 64898 147218 64982 147454
rect 65218 147218 65302 147454
rect 65538 147218 65622 147454
rect 65858 147218 71857 147454
rect 72093 147218 165561 147454
rect 165797 147218 403813 147454
rect 404049 147218 497517 147454
rect 497753 147218 504050 147454
rect 504286 147218 504370 147454
rect 504606 147218 504690 147454
rect 504926 147218 505010 147454
rect 505246 147218 505330 147454
rect 505566 147218 505650 147454
rect 505886 147218 505970 147454
rect 506206 147218 506290 147454
rect 506526 147218 506610 147454
rect 506846 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 63062 147134
rect 63298 146898 63382 147134
rect 63618 146898 63702 147134
rect 63938 146898 64022 147134
rect 64258 146898 64342 147134
rect 64578 146898 64662 147134
rect 64898 146898 64982 147134
rect 65218 146898 65302 147134
rect 65538 146898 65622 147134
rect 65858 146898 71857 147134
rect 72093 146898 165561 147134
rect 165797 146898 403813 147134
rect 404049 146898 497517 147134
rect 497753 146898 504050 147134
rect 504286 146898 504370 147134
rect 504606 146898 504690 147134
rect 504926 146898 505010 147134
rect 505246 146898 505330 147134
rect 505566 146898 505650 147134
rect 505886 146898 505970 147134
rect 506206 146898 506290 147134
rect 506526 146898 506610 147134
rect 506846 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 59062 129454
rect 59298 129218 59382 129454
rect 59618 129218 59702 129454
rect 59938 129218 60022 129454
rect 60258 129218 60342 129454
rect 60578 129218 60662 129454
rect 60898 129218 60982 129454
rect 61218 129218 61302 129454
rect 61538 129218 61622 129454
rect 61858 129218 71177 129454
rect 71413 129218 166241 129454
rect 166477 129218 403133 129454
rect 403369 129218 498197 129454
rect 498433 129218 508050 129454
rect 508286 129218 508370 129454
rect 508606 129218 508690 129454
rect 508926 129218 509010 129454
rect 509246 129218 509330 129454
rect 509566 129218 509650 129454
rect 509886 129218 509970 129454
rect 510206 129218 510290 129454
rect 510526 129218 510610 129454
rect 510846 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 59062 129134
rect 59298 128898 59382 129134
rect 59618 128898 59702 129134
rect 59938 128898 60022 129134
rect 60258 128898 60342 129134
rect 60578 128898 60662 129134
rect 60898 128898 60982 129134
rect 61218 128898 61302 129134
rect 61538 128898 61622 129134
rect 61858 128898 71177 129134
rect 71413 128898 166241 129134
rect 166477 128898 403133 129134
rect 403369 128898 498197 129134
rect 498433 128898 508050 129134
rect 508286 128898 508370 129134
rect 508606 128898 508690 129134
rect 508926 128898 509010 129134
rect 509246 128898 509330 129134
rect 509566 128898 509650 129134
rect 509886 128898 509970 129134
rect 510206 128898 510290 129134
rect 510526 128898 510610 129134
rect 510846 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 63062 111454
rect 63298 111218 63382 111454
rect 63618 111218 63702 111454
rect 63938 111218 64022 111454
rect 64258 111218 64342 111454
rect 64578 111218 64662 111454
rect 64898 111218 64982 111454
rect 65218 111218 65302 111454
rect 65538 111218 65622 111454
rect 65858 111218 71857 111454
rect 72093 111218 165561 111454
rect 165797 111218 403813 111454
rect 404049 111218 497517 111454
rect 497753 111218 504050 111454
rect 504286 111218 504370 111454
rect 504606 111218 504690 111454
rect 504926 111218 505010 111454
rect 505246 111218 505330 111454
rect 505566 111218 505650 111454
rect 505886 111218 505970 111454
rect 506206 111218 506290 111454
rect 506526 111218 506610 111454
rect 506846 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 63062 111134
rect 63298 110898 63382 111134
rect 63618 110898 63702 111134
rect 63938 110898 64022 111134
rect 64258 110898 64342 111134
rect 64578 110898 64662 111134
rect 64898 110898 64982 111134
rect 65218 110898 65302 111134
rect 65538 110898 65622 111134
rect 65858 110898 71857 111134
rect 72093 110898 165561 111134
rect 165797 110898 403813 111134
rect 404049 110898 497517 111134
rect 497753 110898 504050 111134
rect 504286 110898 504370 111134
rect 504606 110898 504690 111134
rect 504926 110898 505010 111134
rect 505246 110898 505330 111134
rect 505566 110898 505650 111134
rect 505886 110898 505970 111134
rect 506206 110898 506290 111134
rect 506526 110898 506610 111134
rect 506846 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 59062 93454
rect 59298 93218 59382 93454
rect 59618 93218 59702 93454
rect 59938 93218 60022 93454
rect 60258 93218 60342 93454
rect 60578 93218 60662 93454
rect 60898 93218 60982 93454
rect 61218 93218 61302 93454
rect 61538 93218 61622 93454
rect 61858 93218 71177 93454
rect 71413 93218 166241 93454
rect 166477 93218 403133 93454
rect 403369 93218 498197 93454
rect 498433 93218 508050 93454
rect 508286 93218 508370 93454
rect 508606 93218 508690 93454
rect 508926 93218 509010 93454
rect 509246 93218 509330 93454
rect 509566 93218 509650 93454
rect 509886 93218 509970 93454
rect 510206 93218 510290 93454
rect 510526 93218 510610 93454
rect 510846 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 59062 93134
rect 59298 92898 59382 93134
rect 59618 92898 59702 93134
rect 59938 92898 60022 93134
rect 60258 92898 60342 93134
rect 60578 92898 60662 93134
rect 60898 92898 60982 93134
rect 61218 92898 61302 93134
rect 61538 92898 61622 93134
rect 61858 92898 71177 93134
rect 71413 92898 166241 93134
rect 166477 92898 403133 93134
rect 403369 92898 498197 93134
rect 498433 92898 508050 93134
rect 508286 92898 508370 93134
rect 508606 92898 508690 93134
rect 508926 92898 509010 93134
rect 509246 92898 509330 93134
rect 509566 92898 509650 93134
rect 509886 92898 509970 93134
rect 510206 92898 510290 93134
rect 510526 92898 510610 93134
rect 510846 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 63062 75454
rect 63298 75218 63382 75454
rect 63618 75218 63702 75454
rect 63938 75218 64022 75454
rect 64258 75218 64342 75454
rect 64578 75218 64662 75454
rect 64898 75218 64982 75454
rect 65218 75218 65302 75454
rect 65538 75218 65622 75454
rect 65858 75218 504050 75454
rect 504286 75218 504370 75454
rect 504606 75218 504690 75454
rect 504926 75218 505010 75454
rect 505246 75218 505330 75454
rect 505566 75218 505650 75454
rect 505886 75218 505970 75454
rect 506206 75218 506290 75454
rect 506526 75218 506610 75454
rect 506846 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 63062 75134
rect 63298 74898 63382 75134
rect 63618 74898 63702 75134
rect 63938 74898 64022 75134
rect 64258 74898 64342 75134
rect 64578 74898 64662 75134
rect 64898 74898 64982 75134
rect 65218 74898 65302 75134
rect 65538 74898 65622 75134
rect 65858 74898 504050 75134
rect 504286 74898 504370 75134
rect 504606 74898 504690 75134
rect 504926 74898 505010 75134
rect 505246 74898 505330 75134
rect 505566 74898 505650 75134
rect 505886 74898 505970 75134
rect 506206 74898 506290 75134
rect 506526 74898 506610 75134
rect 506846 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 59062 57454
rect 59298 57218 59382 57454
rect 59618 57218 59702 57454
rect 59938 57218 60022 57454
rect 60258 57218 60342 57454
rect 60578 57218 60662 57454
rect 60898 57218 60982 57454
rect 61218 57218 61302 57454
rect 61538 57218 61622 57454
rect 61858 57218 508050 57454
rect 508286 57218 508370 57454
rect 508606 57218 508690 57454
rect 508926 57218 509010 57454
rect 509246 57218 509330 57454
rect 509566 57218 509650 57454
rect 509886 57218 509970 57454
rect 510206 57218 510290 57454
rect 510526 57218 510610 57454
rect 510846 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 59062 57134
rect 59298 56898 59382 57134
rect 59618 56898 59702 57134
rect 59938 56898 60022 57134
rect 60258 56898 60342 57134
rect 60578 56898 60662 57134
rect 60898 56898 60982 57134
rect 61218 56898 61302 57134
rect 61538 56898 61622 57134
rect 61858 56898 508050 57134
rect 508286 56898 508370 57134
rect 508606 56898 508690 57134
rect 508926 56898 509010 57134
rect 509246 56898 509330 57134
rect 509566 56898 509650 57134
rect 509886 56898 509970 57134
rect 510206 56898 510290 57134
rect 510526 56898 510610 57134
rect 510846 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 63062 39454
rect 63298 39218 63382 39454
rect 63618 39218 63702 39454
rect 63938 39218 64022 39454
rect 64258 39218 64342 39454
rect 64578 39218 64662 39454
rect 64898 39218 64982 39454
rect 65218 39218 65302 39454
rect 65538 39218 65622 39454
rect 65858 39218 504050 39454
rect 504286 39218 504370 39454
rect 504606 39218 504690 39454
rect 504926 39218 505010 39454
rect 505246 39218 505330 39454
rect 505566 39218 505650 39454
rect 505886 39218 505970 39454
rect 506206 39218 506290 39454
rect 506526 39218 506610 39454
rect 506846 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 63062 39134
rect 63298 38898 63382 39134
rect 63618 38898 63702 39134
rect 63938 38898 64022 39134
rect 64258 38898 64342 39134
rect 64578 38898 64662 39134
rect 64898 38898 64982 39134
rect 65218 38898 65302 39134
rect 65538 38898 65622 39134
rect 65858 38898 504050 39134
rect 504286 38898 504370 39134
rect 504606 38898 504690 39134
rect 504926 38898 505010 39134
rect 505246 38898 505330 39134
rect 505566 38898 505650 39134
rect 505886 38898 505970 39134
rect 506206 38898 506290 39134
rect 506526 38898 506610 39134
rect 506846 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use azadi_soc_top_caravel  mprj
timestamp 0
transform 1 0 55000 0 1 30000
box 0 0 460000 443836
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 475836 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 475836 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 475836 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 475836 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 475836 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 475836 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 475836 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 475836 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 475836 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 475836 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 475836 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 475836 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 475836 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 475836 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 475836 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 475836 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 475836 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 475836 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 475836 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 475836 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 475836 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 475836 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 475836 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 475836 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 475836 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 475836 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 475836 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 475836 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 475836 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 475836 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 475836 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 475836 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 475836 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 475836 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 475836 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 475836 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 475836 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 475836 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 475836 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 475836 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 475836 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 475836 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 475836 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 475836 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 475836 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 475836 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 475836 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 475836 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 475836 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 475836 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 475836 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 475836 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 475836 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 475836 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 475836 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 475836 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 475836 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 475836 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 475836 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 475836 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 475836 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 475836 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 475836 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 475836 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 475836 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 475836 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 475836 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 475836 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 475836 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 475836 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 475836 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 475836 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 475836 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 475836 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 475836 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 475836 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 475836 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 475836 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 475836 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 475836 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 475836 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 475836 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 475836 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 475836 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 475836 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 475836 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 475836 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 475836 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 475836 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 475836 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 475836 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 475836 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 475836 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 475836 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 475836 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 475836 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 475836 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 475836 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 475836 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 475836 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 475836 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 475836 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 475836 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 475836 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
