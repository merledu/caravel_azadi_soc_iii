##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Wed Mar 16 02:15:22 2022
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2300.000000 BY 2219.180000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 241.897 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1291.06 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 4.180000 0.000000 4.320000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.711 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.708 LAYER met2  ;
    ANTENNAMAXAREACAR 26.9062 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.329 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 2.225000 0.000000 2.365000 0.485000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.530000 0.000000 472.670000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.710000 0.000000 158.850000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.120000 0.000000 477.260000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.940000 0.000000 468.080000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.435000 0.000000 463.575000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.930000 0.000000 459.070000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.340000 0.000000 454.480000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.315000 0.000000 304.455000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.640000 0.000000 299.780000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.220000 0.000000 295.360000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.545000 0.000000 290.685000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.125000 0.000000 286.265000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.535000 0.000000 281.675000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.945000 0.000000 277.085000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.440000 0.000000 272.580000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.850000 0.000000 267.990000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.260000 0.000000 263.400000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.840000 0.000000 258.980000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.250000 0.000000 254.390000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.745000 0.000000 249.885000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.155000 0.000000 245.295000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.565000 0.000000 240.705000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.060000 0.000000 236.200000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470000 0.000000 231.610000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.965000 0.000000 227.105000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.460000 0.000000 222.600000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.785000 0.000000 217.925000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.365000 0.000000 213.505000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.690000 0.000000 208.830000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.185000 0.000000 204.325000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.680000 0.000000 199.820000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.175000 0.000000 195.315000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.585000 0.000000 190.725000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.080000 0.000000 186.220000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.405000 0.000000 181.545000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.985000 0.000000 177.125000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.310000 0.000000 172.450000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.890000 0.000000 168.030000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.300000 0.000000 163.440000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.205000 0.000000 154.345000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.615000 0.000000 149.755000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.025000 0.000000 145.165000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.605000 0.000000 140.745000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.015000 0.000000 136.155000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.510000 0.000000 131.650000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.920000 0.000000 127.060000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.330000 0.000000 122.470000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.825000 0.000000 117.965000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.235000 0.000000 113.375000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.730000 0.000000 108.870000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.225000 0.000000 104.365000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.550000 0.000000 99.690000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.215000 0.000000 95.355000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.455000 0.000000 90.595000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.035000 0.000000 86.175000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.445000 0.000000 81.585000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.940000 0.000000 77.080000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.265000 0.000000 72.405000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.845000 0.000000 67.985000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.170000 0.000000 63.310000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.750000 0.000000 58.890000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.075000 0.000000 54.215000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.655000 0.000000 49.795000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.065000 0.000000 45.205000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.560000 0.000000 40.700000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.055000 0.000000 36.195000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.550000 0.000000 31.690000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.960000 0.000000 27.100000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.455000 0.000000 22.595000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.865000 0.000000 18.005000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.275000 0.000000 13.415000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 8.770000 0.000000 8.910000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 449.835000 0.000000 449.975000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 445.160000 0.000000 445.300000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 440.825000 0.000000 440.965000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 436.065000 0.000000 436.205000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 431.645000 0.000000 431.785000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 427.055000 0.000000 427.195000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 422.550000 0.000000 422.690000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 417.960000 0.000000 418.100000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 413.455000 0.000000 413.595000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 408.780000 0.000000 408.920000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 404.360000 0.000000 404.500000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 399.770000 0.000000 399.910000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 395.180000 0.000000 395.320000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 390.675000 0.000000 390.815000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 386.085000 0.000000 386.225000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 381.665000 0.000000 381.805000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 376.990000 0.000000 377.130000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 372.485000 0.000000 372.625000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 367.980000 0.000000 368.120000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 363.390000 0.000000 363.530000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 358.885000 0.000000 359.025000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 354.295000 0.000000 354.435000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 349.705000 0.000000 349.845000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 345.200000 0.000000 345.340000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 340.695000 0.000000 340.835000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 336.020000 0.000000 336.160000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 331.600000 0.000000 331.740000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 326.925000 0.000000 327.065000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 322.590000 0.000000 322.730000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 317.830000 0.000000 317.970000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 313.410000 0.000000 313.550000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 308.820000 0.000000 308.960000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.030000 0.000000 1059.170000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.355000 0.000000 1054.495000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.105000 0.000000 1050.245000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.430000 0.000000 1045.570000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.010000 0.000000 1041.150000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.335000 0.000000 1036.475000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.830000 0.000000 1031.970000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.240000 0.000000 1027.380000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.735000 0.000000 1022.875000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.060000 0.000000 1018.200000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.640000 0.000000 1013.780000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.965000 0.000000 1009.105000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.460000 0.000000 1004.600000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.870000 0.000000 1000.010000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.280000 0.000000 995.420000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.945000 0.000000 991.085000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.355000 0.000000 986.495000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.765000 0.000000 981.905000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.260000 0.000000 977.400000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.670000 0.000000 972.810000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.165000 0.000000 968.305000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.575000 0.000000 963.715000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.985000 0.000000 959.125000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.480000 0.000000 954.620000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.890000 0.000000 950.030000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.300000 0.000000 945.440000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.795000 0.000000 940.935000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.120000 0.000000 936.260000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.870000 0.000000 932.010000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.195000 0.000000 927.335000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.690000 0.000000 922.830000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.100000 0.000000 918.240000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.595000 0.000000 913.735000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.005000 0.000000 909.145000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.500000 0.000000 904.640000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.825000 0.000000 899.965000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.405000 0.000000 895.545000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.730000 0.000000 890.870000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.225000 0.000000 886.365000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.720000 0.000000 881.860000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.045000 0.000000 877.185000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710000 0.000000 872.850000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.120000 0.000000 868.260000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.530000 0.000000 863.670000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.025000 0.000000 859.165000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.435000 0.000000 854.575000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.845000 0.000000 849.985000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.340000 0.000000 845.480000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.750000 0.000000 840.890000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.245000 0.000000 836.385000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.655000 0.000000 831.795000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.065000 0.000000 827.205000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.645000 0.000000 822.785000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.885000 0.000000 818.025000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.635000 0.000000 813.775000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.960000 0.000000 809.100000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.455000 0.000000 804.595000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.865000 0.000000 800.005000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.360000 0.000000 795.500000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.685000 0.000000 790.825000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.265000 0.000000 786.405000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.590000 0.000000 781.730000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.255000 0.000000 777.395000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.495000 0.000000 772.635000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.990000 0.000000 768.130000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.485000 0.000000 763.625000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.810000 0.000000 758.950000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.390000 0.000000 754.530000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.885000 0.000000 750.025000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.295000 0.000000 745.435000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.790000 0.000000 740.930000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.200000 0.000000 736.340000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.610000 0.000000 731.750000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.105000 0.000000 727.245000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.515000 0.000000 722.655000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.925000 0.000000 718.065000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.420000 0.000000 713.560000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.915000 0.000000 709.055000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.410000 0.000000 704.550000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.820000 0.000000 699.960000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.315000 0.000000 695.455000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.725000 0.000000 690.865000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.220000 0.000000 686.360000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.630000 0.000000 681.770000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.125000 0.000000 677.265000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.450000 0.000000 672.590000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.030000 0.000000 668.170000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.355000 0.000000 663.495000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.850000 0.000000 658.990000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.260000 0.000000 654.400000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.840000 0.000000 649.980000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.250000 0.000000 645.390000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.745000 0.000000 640.885000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.155000 0.000000 636.295000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.650000 0.000000 631.790000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.060000 0.000000 627.200000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.555000 0.000000 622.695000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.965000 0.000000 618.105000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.460000 0.000000 613.600000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.870000 0.000000 609.010000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.450000 0.000000 604.590000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.860000 0.000000 600.000000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.355000 0.000000 595.495000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.765000 0.000000 590.905000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.345000 0.000000 586.485000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.670000 0.000000 581.810000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.165000 0.000000 577.305000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.575000 0.000000 572.715000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.070000 0.000000 568.210000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.395000 0.000000 563.535000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.975000 0.000000 559.115000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.300000 0.000000 554.440000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.8835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 25.323 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.379 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 549.965000 0.000000 550.105000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 22.2202 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.802 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 545.290000 0.000000 545.430000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.2175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 15.584 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.7907 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 540.785000 0.000000 540.925000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.6675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 22.7275 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.148 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 536.195000 0.000000 536.335000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.936 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0637 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.0869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.197858 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 531.690000 0.000000 531.830000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.8115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 19.9438 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.5081 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 527.015000 0.000000 527.155000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.7335 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 13.4535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.2985 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 522.595000 0.000000 522.735000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 20.1796 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.3141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 518.005000 0.000000 518.145000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.051 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5834 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.0381 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 513.500000 0.000000 513.640000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.2535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2996 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.1202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 508.910000 0.000000 509.050000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.02 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.884 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4641 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.4417 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 504.320000 0.000000 504.460000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.9835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7598 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.3293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 499.815000 0.000000 499.955000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.8855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 11.426 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.442 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.255272 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 495.225000 0.000000 495.365000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.8925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 20.583 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.7657 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 490.635000 0.000000 490.775000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.7215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.9863 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.7832 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 486.215000 0.000000 486.355000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.2025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 13.3821 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.9469 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 481.625000 0.000000 481.765000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1641.110000 0.000000 1641.250000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1636.520000 0.000000 1636.660000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1632.015000 0.000000 1632.155000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1627.340000 0.000000 1627.480000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1622.920000 0.000000 1623.060000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1618.245000 0.000000 1618.385000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1613.910000 0.000000 1614.050000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1609.235000 0.000000 1609.375000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1604.730000 0.000000 1604.870000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1600.140000 0.000000 1600.280000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1595.550000 0.000000 1595.690000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1591.045000 0.000000 1591.185000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1586.455000 0.000000 1586.595000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1581.950000 0.000000 1582.090000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1577.445000 0.000000 1577.585000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1572.855000 0.000000 1572.995000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1568.265000 0.000000 1568.405000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1563.845000 0.000000 1563.985000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1559.170000 0.000000 1559.310000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1554.750000 0.000000 1554.890000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1550.160000 0.000000 1550.300000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1545.570000 0.000000 1545.710000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1541.065000 0.000000 1541.205000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1536.390000 0.000000 1536.530000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1531.885000 0.000000 1532.025000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1527.295000 0.000000 1527.435000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1522.875000 0.000000 1523.015000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1518.285000 0.000000 1518.425000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1513.780000 0.000000 1513.920000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1509.105000 0.000000 1509.245000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1504.770000 0.000000 1504.910000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1500.010000 0.000000 1500.150000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1495.675000 0.000000 1495.815000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1491.000000 0.000000 1491.140000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1486.495000 0.000000 1486.635000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1481.905000 0.000000 1482.045000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1477.315000 0.000000 1477.455000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1472.725000 0.000000 1472.865000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1468.220000 0.000000 1468.360000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1463.715000 0.000000 1463.855000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1459.210000 0.000000 1459.350000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1454.620000 0.000000 1454.760000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1450.030000 0.000000 1450.170000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1445.610000 0.000000 1445.750000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1440.935000 0.000000 1441.075000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1436.430000 0.000000 1436.570000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1431.925000 0.000000 1432.065000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1427.335000 0.000000 1427.475000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1422.830000 0.000000 1422.970000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1418.155000 0.000000 1418.295000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1413.650000 0.000000 1413.790000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1409.060000 0.000000 1409.200000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1404.640000 0.000000 1404.780000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1399.965000 0.000000 1400.105000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1395.545000 0.000000 1395.685000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1390.870000 0.000000 1391.010000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1386.535000 0.000000 1386.675000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1381.775000 0.000000 1381.915000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1377.355000 0.000000 1377.495000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1372.765000 0.000000 1372.905000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1368.260000 0.000000 1368.400000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1363.670000 0.000000 1363.810000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1359.080000 0.000000 1359.220000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1354.490000 0.000000 1354.630000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1349.985000 0.000000 1350.125000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1345.480000 0.000000 1345.620000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1340.890000 0.000000 1341.030000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1336.385000 0.000000 1336.525000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1331.795000 0.000000 1331.935000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1327.375000 0.000000 1327.515000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1322.785000 0.000000 1322.925000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1318.195000 0.000000 1318.335000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1313.690000 0.000000 1313.830000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1309.100000 0.000000 1309.240000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1304.510000 0.000000 1304.650000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1299.920000 0.000000 1300.060000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1295.415000 0.000000 1295.555000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1290.825000 0.000000 1290.965000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1286.405000 0.000000 1286.545000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1281.730000 0.000000 1281.870000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1277.310000 0.000000 1277.450000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1272.635000 0.000000 1272.775000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1268.300000 0.000000 1268.440000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1263.625000 0.000000 1263.765000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1259.120000 0.000000 1259.260000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1254.530000 0.000000 1254.670000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1250.025000 0.000000 1250.165000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1245.350000 0.000000 1245.490000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1240.845000 0.000000 1240.985000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1236.255000 0.000000 1236.395000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1231.750000 0.000000 1231.890000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1227.245000 0.000000 1227.385000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1222.655000 0.000000 1222.795000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1218.235000 0.000000 1218.375000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1213.560000 0.000000 1213.700000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1208.970000 0.000000 1209.110000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1204.550000 0.000000 1204.690000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1199.960000 0.000000 1200.100000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1195.455000 0.000000 1195.595000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1190.865000 0.000000 1191.005000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1186.360000 0.000000 1186.500000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1181.770000 0.000000 1181.910000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1177.265000 0.000000 1177.405000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1172.590000 0.000000 1172.730000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1168.340000 0.000000 1168.480000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1163.580000 0.000000 1163.720000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1159.245000 0.000000 1159.385000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1154.570000 0.000000 1154.710000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1150.065000 0.000000 1150.205000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1145.475000 0.000000 1145.615000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1140.970000 0.000000 1141.110000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1136.380000 0.000000 1136.520000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1131.875000 0.000000 1132.015000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1127.200000 0.000000 1127.340000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1122.695000 0.000000 1122.835000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1118.105000 0.000000 1118.245000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1113.515000 0.000000 1113.655000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1109.180000 0.000000 1109.320000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1104.505000 0.000000 1104.645000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1100.085000 0.000000 1100.225000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1095.495000 0.000000 1095.635000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1090.905000 0.000000 1091.045000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1086.400000 0.000000 1086.540000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1081.810000 0.000000 1081.950000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1077.220000 0.000000 1077.360000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1072.715000 0.000000 1072.855000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.516 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.24 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1068.125000 0.000000 1068.265000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1063.535000 0.000000 1063.675000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2223.190000 0.000000 2223.330000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.515000 0.000000 2218.655000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.010000 0.000000 2214.150000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.420000 0.000000 2209.560000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.915000 0.000000 2205.055000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2200.325000 0.000000 2200.465000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.735000 0.000000 2195.875000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.145000 0.000000 2191.285000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.640000 0.000000 2186.780000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2182.050000 0.000000 2182.190000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.630000 0.000000 2177.770000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.125000 0.000000 2173.265000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.450000 0.000000 2168.590000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.030000 0.000000 2164.170000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.440000 0.000000 2159.580000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.850000 0.000000 2154.990000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2150.345000 0.000000 2150.485000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.755000 0.000000 2145.895000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.250000 0.000000 2141.390000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.575000 0.000000 2136.715000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2132.070000 0.000000 2132.210000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2127.480000 0.000000 2127.620000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.975000 0.000000 2123.115000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.300000 0.000000 2118.440000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2114.050000 0.000000 2114.190000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.375000 0.000000 2109.515000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.955000 0.000000 2105.095000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.280000 0.000000 2100.420000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.775000 0.000000 2095.915000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.185000 0.000000 2091.325000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.680000 0.000000 2086.820000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.005000 0.000000 2082.145000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.500000 0.000000 2077.640000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.910000 0.000000 2073.050000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.405000 0.000000 2068.545000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.815000 0.000000 2063.955000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.140000 0.000000 2059.280000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.890000 0.000000 2055.030000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2050.300000 0.000000 2050.440000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.795000 0.000000 2045.935000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.205000 0.000000 2041.345000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.615000 0.000000 2036.755000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2032.110000 0.000000 2032.250000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.520000 0.000000 2027.660000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.930000 0.000000 2023.070000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.340000 0.000000 2018.480000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.835000 0.000000 2013.975000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.245000 0.000000 2009.385000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.825000 0.000000 2004.965000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.065000 0.000000 2000.205000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.815000 0.000000 1995.955000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.140000 0.000000 1991.280000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.635000 0.000000 1986.775000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.045000 0.000000 1982.185000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.540000 0.000000 1977.680000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.950000 0.000000 1973.090000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.445000 0.000000 1968.585000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.770000 0.000000 1963.910000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.265000 0.000000 1959.405000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.675000 0.000000 1954.815000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.170000 0.000000 1950.310000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.665000 0.000000 1945.805000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.905000 0.000000 1941.045000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.655000 0.000000 1936.795000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.065000 0.000000 1932.205000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.475000 0.000000 1927.615000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.970000 0.000000 1923.110000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.380000 0.000000 1918.520000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.875000 0.000000 1914.015000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.285000 0.000000 1909.425000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.695000 0.000000 1904.835000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.105000 0.000000 1900.245000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.600000 0.000000 1895.740000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.925000 0.000000 1891.065000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.590000 0.000000 1886.730000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.830000 0.000000 1881.970000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.580000 0.000000 1877.720000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.905000 0.000000 1873.045000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.400000 0.000000 1868.540000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.810000 0.000000 1863.950000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.305000 0.000000 1859.445000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.630000 0.000000 1854.770000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.210000 0.000000 1850.350000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.535000 0.000000 1845.675000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.030000 0.000000 1841.170000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.440000 0.000000 1836.580000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.765000 0.000000 1831.905000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.430000 0.000000 1827.570000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.670000 0.000000 1822.810000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.420000 0.000000 1818.560000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.830000 0.000000 1813.970000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.240000 0.000000 1809.380000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.735000 0.000000 1804.875000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.145000 0.000000 1800.285000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.555000 0.000000 1795.695000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.050000 0.000000 1791.190000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.460000 0.000000 1786.600000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.870000 0.000000 1782.010000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.365000 0.000000 1777.505000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.860000 0.000000 1773.000000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.355000 0.000000 1768.495000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.765000 0.000000 1763.905000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1759.345000 0.000000 1759.485000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.755000 0.000000 1754.895000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.250000 0.000000 1750.390000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.660000 0.000000 1745.800000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.155000 0.000000 1741.295000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.480000 0.000000 1736.620000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.145000 0.000000 1732.285000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.385000 0.000000 1727.525000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.965000 0.000000 1723.105000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.375000 0.000000 1718.515000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.785000 0.000000 1713.925000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.280000 0.000000 1709.420000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.690000 0.000000 1704.830000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.185000 0.000000 1700.325000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.680000 0.000000 1695.820000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.090000 0.000000 1691.230000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.585000 0.000000 1686.725000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.995000 0.000000 1682.135000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.405000 0.000000 1677.545000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.985000 0.000000 1673.125000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.395000 0.000000 1668.535000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.805000 0.000000 1663.945000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1659.300000 0.000000 1659.440000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.625000 0.000000 1654.765000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.205000 0.000000 1650.345000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.530000 0.000000 1645.670000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 57.420000 0.800000 57.720000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.0074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 187.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.3668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 391.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 111.392 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 570.545 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.532248 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 205.150000 0.800000 205.450000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 143.787 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 769.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 211.56 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1095.8 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.673088 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 328.450000 0.800000 328.750000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9066 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 97.9572 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 526.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 128.817 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 668.836 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.532248 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 492.850000 0.800000 493.150000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 314.901 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1679.94 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.2816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 125.419 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 652.958 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.599775 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 657.250000 0.800000 657.550000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225.376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1203.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.9432 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 36.3992 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 164.078 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.494517 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 821.650000 0.800000 821.950000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 253.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1352.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.1304 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 73.5627 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.494517 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 985.950000 0.800000 986.250000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.1406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 283.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.7712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 427.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 131.598 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 670.264 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.682086 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1150.450000 0.800000 1150.750000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 68.7438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 367.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 102.183 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 532.298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.494517 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1314.750000 0.800000 1315.050000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.2092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 220.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 34.8985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 158.124 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1479.150000 0.800000 1479.450000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.4824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.765 LAYER met3  ;
    ANTENNAMAXAREACAR 98.8391 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 473.61 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.670057 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.5158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.888 LAYER met4  ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 150.263 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 748.38 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1643.550000 0.800000 1643.850000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1807.950000 0.800000 1808.250000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6513 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 62.4012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 334.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 115.531 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 610.14 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.19028 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1972.350000 0.800000 1972.650000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 69.0456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 369.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 156.831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 823.003 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2136.650000 0.800000 2136.950000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 111.934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 559.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 57.9546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 310.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 147.111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 761.589 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 127.855000 2218.690000 127.995000 2219.180000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 110.837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 553.906 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 65.3454 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 349.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 93.9968 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 489.996 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 383.960000 2218.690000 384.100000 2219.180000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 116.862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 584.031 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 56.5626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 302.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 113.646 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 572.066 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.14743 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 640.235000 2218.690000 640.375000 2219.180000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 115.889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 579.166 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 56.4186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 101.338 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 509.508 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 896.595000 2218.690000 896.735000 2219.180000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 115.981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 579.743 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.2048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.765 LAYER met3  ;
    ANTENNAMAXAREACAR 54.1069 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 252.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.921942 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.7418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 361.76 LAYER met4  ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 127.421 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 643.779 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.921942 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1152.700000 2218.690000 1152.840000 2219.180000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 106.111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 530.274 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.709 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.9794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 363.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 135.147 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 706.38 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.46806 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1408.890000 2218.690000 1409.030000 2219.180000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 91.2142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 455.91 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 90.385 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 482.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.7816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 479.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 150.421 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 782.232 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1665.165000 2218.690000 1665.305000 2219.180000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 537.957 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 68.2746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 365.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 99.189 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 496.763 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1921.355000 2218.690000 1921.495000 2219.180000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 110.68 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 553.122 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.6018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 342.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 91.2335 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 480.005 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.46806 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2177.630000 2218.690000 2177.770000 2219.180000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 68.448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 367.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 116.196 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 598.684 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.46806 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 2094.050000 2300.000000 2094.350000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0203 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 83.075 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 428.128 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04451 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1926.450000 2300.000000 1926.750000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7967 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met3  ;
    ANTENNAMAXAREACAR 112.414 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 540.569 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.691083 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1758.950000 2300.000000 1759.250000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.0322 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met3  ;
    ANTENNAMAXAREACAR 74.2435 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.28 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1591.350000 2300.000000 1591.650000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 68.0164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 363.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 66.5715 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 358.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 97.1644 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 504.564 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1423.750000 2300.000000 1424.050000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 88.3402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 472.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 22.5716 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 88.1513 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.443525 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1256.350000 2300.000000 1256.650000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 226.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1210.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 57.3359 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.247 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.673088 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1088.750000 2300.000000 1089.050000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 40.7634 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.659 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 921.250000 2300.000000 921.550000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 753.650000 2300.000000 753.950000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 69.0395 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 368.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.7388 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 149.438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 799.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 715.404 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 3722.11 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 627.950000 2300.000000 628.250000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 502.350000 2300.000000 502.650000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met3  ;
    ANTENNAMAXAREACAR 39.6031 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.194 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 376.650000 2300.000000 376.950000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.8334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.2228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 91.6404 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 452.743 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 250.950000 2300.000000 251.250000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.4314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met4  ;
    ANTENNAMAXAREACAR 39.0249 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.623 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.599775 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 125.350000 2300.000000 125.650000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 3.950000 2300.000000 4.250000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 40.850000 0.800000 41.150000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.050000 0.800000 164.350000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.1352 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 287.450000 0.800000 287.750000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 451.750000 0.800000 452.050000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.9036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 616.150000 0.800000 616.450000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 268.359 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1431.71 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.7286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.16 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 780.450000 0.800000 780.750000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 255.839 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1365.41 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.9916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 304.896 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 944.950000 0.800000 945.250000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 156.24 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 833.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.2314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.312 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1109.250000 0.800000 1109.550000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.1542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 193.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1273.750000 0.800000 1274.050000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 98.3208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 524.848 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1438.050000 0.800000 1438.350000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1602.450000 0.800000 1602.750000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1766.850000 0.800000 1767.150000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1931.150000 0.800000 1931.450000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.5504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2095.650000 0.800000 2095.950000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 70.6803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 353.294 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.765000 2218.690000 63.905000 2219.180000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.7765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 319.955000 2218.690000 320.095000 2219.180000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 118.672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 593.079 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.6598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 576.145000 2218.690000 576.285000 2219.180000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 50.329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 251.419 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 832.420000 2218.690000 832.560000 2219.180000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 32.8186 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 163.513 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1088.610000 2218.690000 1088.750000 2219.180000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 108.199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 540.834 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.9768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 405.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3915 LAYER met4  ;
    ANTENNAMAXAREACAR 236.728 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1252.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.561287 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1344.885000 2218.690000 1345.025000 2219.180000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 86.3758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 431.718 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.575 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.2808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1601.075000 2218.690000 1601.215000 2219.180000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.6536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 98.042 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1857.350000 2218.690000 1857.490000 2219.180000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.5279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.4135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2113.455000 2218.690000 2113.595000 2219.180000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 2135.950000 2300.000000 2136.250000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.7172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 313.624 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1968.450000 2300.000000 1968.750000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1800.750000 2300.000000 1801.050000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1633.250000 2300.000000 1633.550000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 82.2372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 439.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1465.750000 2300.000000 1466.050000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 141.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 753.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1298.150000 2300.000000 1298.450000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.84 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1130.650000 2300.000000 1130.950000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 963.150000 2300.000000 963.450000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 795.550000 2300.000000 795.850000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 669.950000 2300.000000 670.250000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.813 LAYER met3  ;
    ANTENNAMAXAREACAR 79.8086 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 391.174 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.555463 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 544.250000 2300.000000 544.550000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8142 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 418.550000 2300.000000 418.850000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 292.950000 2300.000000 293.250000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 167.250000 2300.000000 167.550000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 41.650000 2300.000000 41.950000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2.150000 0.800000 2.450000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 61.0974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 325.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 123.050000 0.800000 123.350000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 246.350000 0.800000 246.650000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 79.2064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 422.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.1334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.456 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 410.650000 0.800000 410.950000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.5026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.5006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.944 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 575.150000 0.800000 575.450000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 739.450000 0.800000 739.750000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.0332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 903.850000 0.800000 904.150000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 149.844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 799.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1068.250000 0.800000 1068.550000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.9278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.752 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1232.550000 0.800000 1232.850000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1396.950000 0.800000 1397.250000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.0578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 374.112 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1561.350000 0.800000 1561.650000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1725.750000 0.800000 1726.050000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1890.150000 0.800000 1890.450000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.9314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2054.450000 0.800000 2054.750000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.394 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.540000 2218.695000 5.680000 2219.180000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.9709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.7465 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 255.865000 2218.690000 256.005000 2219.180000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.9235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 512.055000 2218.690000 512.195000 2219.180000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 111.85 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 558.905 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 768.245000 2218.690000 768.385000 2219.180000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 65.284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 326.312 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1024.520000 2218.690000 1024.660000 2219.180000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 105.675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 528.15 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1280.710000 2218.690000 1280.850000 2219.180000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 91.1292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 455.42 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1537.070000 2218.690000 1537.210000 2219.180000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 92.3347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 461.395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1793.260000 2218.690000 1793.400000 2219.180000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.0717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.2505 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2049.365000 2218.690000 2049.505000 2219.180000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6626 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.6734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 2176.150000 2300.000000 2176.450000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.2574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 2010.250000 2300.000000 2010.550000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.6654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1842.750000 2300.000000 1843.050000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1675.150000 2300.000000 1675.450000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.304 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1507.550000 2300.000000 1507.850000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1340.050000 2300.000000 1340.350000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1172.550000 2300.000000 1172.850000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.56 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1004.950000 2300.000000 1005.250000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 837.450000 2300.000000 837.750000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.56 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 711.750000 2300.000000 712.050000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 586.150000 2300.000000 586.450000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 460.450000 2300.000000 460.750000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 334.750000 2300.000000 335.050000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.8124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 212.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 209.150000 2300.000000 209.450000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0036 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 83.550000 2300.000000 83.850000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 369.550000 0.800000 369.850000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 533.950000 0.800000 534.250000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 698.350000 0.800000 698.650000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 862.750000 0.800000 863.050000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1027.150000 0.800000 1027.450000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1191.550000 0.800000 1191.850000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1355.850000 0.800000 1356.150000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1520.350000 0.800000 1520.650000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1684.550000 0.800000 1684.850000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1849.050000 0.800000 1849.350000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2013.350000 0.800000 2013.650000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2175.750000 0.800000 2176.050000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.775000 2218.690000 191.915000 2219.180000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.220000 2218.690000 448.360000 2219.180000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.155000 2218.690000 704.295000 2219.180000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.515000 2218.690000 960.655000 2219.180000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.620000 2218.690000 1216.760000 2219.180000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.895000 2218.690000 1473.035000 2219.180000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.085000 2218.690000 1729.225000 2219.180000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.445000 2218.690000 1985.585000 2219.180000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.405000 2218.695000 2238.545000 2219.180000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 2052.150000 2300.000000 2052.450000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1884.550000 2300.000000 1884.850000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1717.050000 2300.000000 1717.350000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1549.450000 2300.000000 1549.750000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1381.950000 2300.000000 1382.250000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1214.350000 2300.000000 1214.650000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 1046.950000 2300.000000 1047.250000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2299.200000 879.350000 2300.000000 879.650000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2227.525000 0.000000 2227.665000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2239.425000 0.000000 2239.565000 0.485000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1750.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2236.620000 0.000000 2236.760000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 350.496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1749.99 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2232.285000 0.000000 2232.425000 0.490000 ;
    END
  END user_irq[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2264.740000 19.840000 2279.740000 2196.960000 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.800000 19.840000 34.800000 2196.960000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2215.705000 234.870000 2217.445000 629.650000 ;
      LAYER met3 ;
        RECT 1740.385000 234.870000 2217.445000 236.610000 ;
      LAYER met3 ;
        RECT 1740.385000 627.910000 2217.445000 629.650000 ;
      LAYER met4 ;
        RECT 1740.385000 234.870000 1742.125000 629.650000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2215.705000 732.370000 2217.445000 1127.150000 ;
      LAYER met3 ;
        RECT 1740.385000 732.370000 2217.445000 734.110000 ;
      LAYER met3 ;
        RECT 1740.385000 1125.410000 2217.445000 1127.150000 ;
      LAYER met4 ;
        RECT 1740.385000 732.370000 1742.125000 1127.150000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2215.705000 1229.870000 2217.445000 1624.650000 ;
      LAYER met3 ;
        RECT 1740.385000 1229.870000 2217.445000 1231.610000 ;
      LAYER met3 ;
        RECT 1740.385000 1622.910000 2217.445000 1624.650000 ;
      LAYER met4 ;
        RECT 1740.385000 1229.870000 1742.125000 1624.650000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2215.705000 1727.370000 2217.445000 2122.150000 ;
      LAYER met3 ;
        RECT 1740.385000 1727.370000 2217.445000 1729.110000 ;
      LAYER met3 ;
        RECT 1740.385000 2120.410000 2217.445000 2122.150000 ;
      LAYER met4 ;
        RECT 1740.385000 1727.370000 1742.125000 2122.150000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 555.925000 234.870000 557.665000 629.650000 ;
      LAYER met3 ;
        RECT 80.605000 234.870000 557.665000 236.610000 ;
      LAYER met3 ;
        RECT 80.605000 627.910000 557.665000 629.650000 ;
      LAYER met4 ;
        RECT 80.605000 234.870000 82.345000 629.650000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 555.925000 732.370000 557.665000 1127.150000 ;
      LAYER met3 ;
        RECT 80.605000 732.370000 557.665000 734.110000 ;
      LAYER met3 ;
        RECT 80.605000 1125.410000 557.665000 1127.150000 ;
      LAYER met4 ;
        RECT 80.605000 732.370000 82.345000 1127.150000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 555.925000 1229.870000 557.665000 1624.650000 ;
      LAYER met3 ;
        RECT 80.605000 1229.870000 557.665000 1231.610000 ;
      LAYER met3 ;
        RECT 80.605000 1622.910000 557.665000 1624.650000 ;
      LAYER met4 ;
        RECT 80.605000 1229.870000 82.345000 1624.650000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 555.925000 1727.370000 557.665000 2122.150000 ;
      LAYER met3 ;
        RECT 80.605000 1727.370000 557.665000 1729.110000 ;
      LAYER met3 ;
        RECT 80.605000 2120.410000 557.665000 2122.150000 ;
      LAYER met4 ;
        RECT 80.605000 1727.370000 82.345000 2122.150000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2244.740000 39.840000 2259.740000 2176.960000 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.800000 39.840000 54.800000 2176.960000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1743.785000 624.510000 2214.045000 626.250000 ;
      LAYER met3 ;
        RECT 1743.785000 238.270000 2214.045000 240.010000 ;
      LAYER met4 ;
        RECT 1743.785000 238.270000 1745.525000 626.250000 ;
      LAYER met4 ;
        RECT 2212.305000 238.270000 2214.045000 626.250000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1743.785000 1122.010000 2214.045000 1123.750000 ;
      LAYER met3 ;
        RECT 1743.785000 735.770000 2214.045000 737.510000 ;
      LAYER met4 ;
        RECT 1743.785000 735.770000 1745.525000 1123.750000 ;
      LAYER met4 ;
        RECT 2212.305000 735.770000 2214.045000 1123.750000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1743.785000 1619.510000 2214.045000 1621.250000 ;
      LAYER met3 ;
        RECT 1743.785000 1233.270000 2214.045000 1235.010000 ;
      LAYER met4 ;
        RECT 1743.785000 1233.270000 1745.525000 1621.250000 ;
      LAYER met4 ;
        RECT 2212.305000 1233.270000 2214.045000 1621.250000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1743.785000 2117.010000 2214.045000 2118.750000 ;
      LAYER met3 ;
        RECT 1743.785000 1730.770000 2214.045000 1732.510000 ;
      LAYER met4 ;
        RECT 1743.785000 1730.770000 1745.525000 2118.750000 ;
      LAYER met4 ;
        RECT 2212.305000 1730.770000 2214.045000 2118.750000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 84.005000 624.510000 554.265000 626.250000 ;
      LAYER met3 ;
        RECT 84.005000 238.270000 554.265000 240.010000 ;
      LAYER met4 ;
        RECT 84.005000 238.270000 85.745000 626.250000 ;
      LAYER met4 ;
        RECT 552.525000 238.270000 554.265000 626.250000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 84.005000 1122.010000 554.265000 1123.750000 ;
      LAYER met3 ;
        RECT 84.005000 735.770000 554.265000 737.510000 ;
      LAYER met4 ;
        RECT 84.005000 735.770000 85.745000 1123.750000 ;
      LAYER met4 ;
        RECT 552.525000 735.770000 554.265000 1123.750000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 84.005000 1619.510000 554.265000 1621.250000 ;
      LAYER met3 ;
        RECT 84.005000 1233.270000 554.265000 1235.010000 ;
      LAYER met4 ;
        RECT 84.005000 1233.270000 85.745000 1621.250000 ;
      LAYER met4 ;
        RECT 552.525000 1233.270000 554.265000 1621.250000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 84.005000 2117.010000 554.265000 2118.750000 ;
      LAYER met3 ;
        RECT 84.005000 1730.770000 554.265000 1732.510000 ;
      LAYER met4 ;
        RECT 84.005000 1730.770000 85.745000 2118.750000 ;
      LAYER met4 ;
        RECT 552.525000 1730.770000 554.265000 2118.750000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2300.000000 2219.180000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2300.000000 2219.180000 ;
    LAYER met2 ;
      RECT 2238.685000 2218.555000 2300.000000 2219.180000 ;
      RECT 2177.910000 2218.555000 2238.265000 2219.180000 ;
      RECT 5.820000 2218.555000 63.625000 2219.180000 ;
      RECT 0.000000 2218.555000 5.400000 2219.180000 ;
      RECT 2177.910000 2218.550000 2300.000000 2218.555000 ;
      RECT 2113.735000 2218.550000 2177.490000 2219.180000 ;
      RECT 2049.645000 2218.550000 2113.315000 2219.180000 ;
      RECT 1985.725000 2218.550000 2049.225000 2219.180000 ;
      RECT 1921.635000 2218.550000 1985.305000 2219.180000 ;
      RECT 1857.630000 2218.550000 1921.215000 2219.180000 ;
      RECT 1793.540000 2218.550000 1857.210000 2219.180000 ;
      RECT 1729.365000 2218.550000 1793.120000 2219.180000 ;
      RECT 1665.445000 2218.550000 1728.945000 2219.180000 ;
      RECT 1601.355000 2218.550000 1665.025000 2219.180000 ;
      RECT 1537.350000 2218.550000 1600.935000 2219.180000 ;
      RECT 1473.175000 2218.550000 1536.930000 2219.180000 ;
      RECT 1409.170000 2218.550000 1472.755000 2219.180000 ;
      RECT 1345.165000 2218.550000 1408.750000 2219.180000 ;
      RECT 1280.990000 2218.550000 1344.745000 2219.180000 ;
      RECT 1216.900000 2218.550000 1280.570000 2219.180000 ;
      RECT 1152.980000 2218.550000 1216.480000 2219.180000 ;
      RECT 1088.890000 2218.550000 1152.560000 2219.180000 ;
      RECT 1024.800000 2218.550000 1088.470000 2219.180000 ;
      RECT 960.795000 2218.550000 1024.380000 2219.180000 ;
      RECT 896.875000 2218.550000 960.375000 2219.180000 ;
      RECT 832.700000 2218.550000 896.455000 2219.180000 ;
      RECT 768.525000 2218.550000 832.280000 2219.180000 ;
      RECT 704.435000 2218.550000 768.105000 2219.180000 ;
      RECT 640.515000 2218.550000 704.015000 2219.180000 ;
      RECT 576.425000 2218.550000 640.095000 2219.180000 ;
      RECT 512.335000 2218.550000 576.005000 2219.180000 ;
      RECT 448.500000 2218.550000 511.915000 2219.180000 ;
      RECT 384.240000 2218.550000 448.080000 2219.180000 ;
      RECT 320.235000 2218.550000 383.820000 2219.180000 ;
      RECT 256.145000 2218.550000 319.815000 2219.180000 ;
      RECT 192.055000 2218.550000 255.725000 2219.180000 ;
      RECT 128.135000 2218.550000 191.635000 2219.180000 ;
      RECT 64.045000 2218.550000 127.715000 2219.180000 ;
      RECT 0.000000 2218.550000 63.625000 2218.555000 ;
      RECT 0.000000 0.630000 2300.000000 2218.550000 ;
      RECT 2236.900000 0.625000 2300.000000 0.630000 ;
      RECT 0.000000 0.625000 4.040000 0.630000 ;
      RECT 2239.705000 0.000000 2300.000000 0.625000 ;
      RECT 2236.900000 0.000000 2239.285000 0.625000 ;
      RECT 2232.565000 0.000000 2236.480000 0.630000 ;
      RECT 2227.805000 0.000000 2232.145000 0.630000 ;
      RECT 2223.470000 0.000000 2227.385000 0.630000 ;
      RECT 2218.795000 0.000000 2223.050000 0.630000 ;
      RECT 2214.290000 0.000000 2218.375000 0.630000 ;
      RECT 2209.700000 0.000000 2213.870000 0.630000 ;
      RECT 2205.195000 0.000000 2209.280000 0.630000 ;
      RECT 2200.605000 0.000000 2204.775000 0.630000 ;
      RECT 2196.015000 0.000000 2200.185000 0.630000 ;
      RECT 2191.425000 0.000000 2195.595000 0.630000 ;
      RECT 2186.920000 0.000000 2191.005000 0.630000 ;
      RECT 2182.330000 0.000000 2186.500000 0.630000 ;
      RECT 2177.910000 0.000000 2181.910000 0.630000 ;
      RECT 2173.405000 0.000000 2177.490000 0.630000 ;
      RECT 2168.730000 0.000000 2172.985000 0.630000 ;
      RECT 2164.310000 0.000000 2168.310000 0.630000 ;
      RECT 2159.720000 0.000000 2163.890000 0.630000 ;
      RECT 2155.130000 0.000000 2159.300000 0.630000 ;
      RECT 2150.625000 0.000000 2154.710000 0.630000 ;
      RECT 2146.035000 0.000000 2150.205000 0.630000 ;
      RECT 2141.530000 0.000000 2145.615000 0.630000 ;
      RECT 2136.855000 0.000000 2141.110000 0.630000 ;
      RECT 2132.350000 0.000000 2136.435000 0.630000 ;
      RECT 2127.760000 0.000000 2131.930000 0.630000 ;
      RECT 2123.255000 0.000000 2127.340000 0.630000 ;
      RECT 2118.580000 0.000000 2122.835000 0.630000 ;
      RECT 2114.330000 0.000000 2118.160000 0.630000 ;
      RECT 2109.655000 0.000000 2113.910000 0.630000 ;
      RECT 2105.235000 0.000000 2109.235000 0.630000 ;
      RECT 2100.560000 0.000000 2104.815000 0.630000 ;
      RECT 2096.055000 0.000000 2100.140000 0.630000 ;
      RECT 2091.465000 0.000000 2095.635000 0.630000 ;
      RECT 2086.960000 0.000000 2091.045000 0.630000 ;
      RECT 2082.285000 0.000000 2086.540000 0.630000 ;
      RECT 2077.780000 0.000000 2081.865000 0.630000 ;
      RECT 2073.190000 0.000000 2077.360000 0.630000 ;
      RECT 2068.685000 0.000000 2072.770000 0.630000 ;
      RECT 2064.095000 0.000000 2068.265000 0.630000 ;
      RECT 2059.420000 0.000000 2063.675000 0.630000 ;
      RECT 2055.170000 0.000000 2059.000000 0.630000 ;
      RECT 2050.580000 0.000000 2054.750000 0.630000 ;
      RECT 2046.075000 0.000000 2050.160000 0.630000 ;
      RECT 2041.485000 0.000000 2045.655000 0.630000 ;
      RECT 2036.895000 0.000000 2041.065000 0.630000 ;
      RECT 2032.390000 0.000000 2036.475000 0.630000 ;
      RECT 2027.800000 0.000000 2031.970000 0.630000 ;
      RECT 2023.210000 0.000000 2027.380000 0.630000 ;
      RECT 2018.620000 0.000000 2022.790000 0.630000 ;
      RECT 2014.115000 0.000000 2018.200000 0.630000 ;
      RECT 2009.525000 0.000000 2013.695000 0.630000 ;
      RECT 2005.105000 0.000000 2009.105000 0.630000 ;
      RECT 2000.345000 0.000000 2004.685000 0.630000 ;
      RECT 1996.095000 0.000000 1999.925000 0.630000 ;
      RECT 1991.420000 0.000000 1995.675000 0.630000 ;
      RECT 1986.915000 0.000000 1991.000000 0.630000 ;
      RECT 1982.325000 0.000000 1986.495000 0.630000 ;
      RECT 1977.820000 0.000000 1981.905000 0.630000 ;
      RECT 1973.230000 0.000000 1977.400000 0.630000 ;
      RECT 1968.725000 0.000000 1972.810000 0.630000 ;
      RECT 1964.050000 0.000000 1968.305000 0.630000 ;
      RECT 1959.545000 0.000000 1963.630000 0.630000 ;
      RECT 1954.955000 0.000000 1959.125000 0.630000 ;
      RECT 1950.450000 0.000000 1954.535000 0.630000 ;
      RECT 1945.945000 0.000000 1950.030000 0.630000 ;
      RECT 1941.185000 0.000000 1945.525000 0.630000 ;
      RECT 1936.935000 0.000000 1940.765000 0.630000 ;
      RECT 1932.345000 0.000000 1936.515000 0.630000 ;
      RECT 1927.755000 0.000000 1931.925000 0.630000 ;
      RECT 1923.250000 0.000000 1927.335000 0.630000 ;
      RECT 1918.660000 0.000000 1922.830000 0.630000 ;
      RECT 1914.155000 0.000000 1918.240000 0.630000 ;
      RECT 1909.565000 0.000000 1913.735000 0.630000 ;
      RECT 1904.975000 0.000000 1909.145000 0.630000 ;
      RECT 1900.385000 0.000000 1904.555000 0.630000 ;
      RECT 1895.880000 0.000000 1899.965000 0.630000 ;
      RECT 1891.205000 0.000000 1895.460000 0.630000 ;
      RECT 1886.870000 0.000000 1890.785000 0.630000 ;
      RECT 1882.110000 0.000000 1886.450000 0.630000 ;
      RECT 1877.860000 0.000000 1881.690000 0.630000 ;
      RECT 1873.185000 0.000000 1877.440000 0.630000 ;
      RECT 1868.680000 0.000000 1872.765000 0.630000 ;
      RECT 1864.090000 0.000000 1868.260000 0.630000 ;
      RECT 1859.585000 0.000000 1863.670000 0.630000 ;
      RECT 1854.910000 0.000000 1859.165000 0.630000 ;
      RECT 1850.490000 0.000000 1854.490000 0.630000 ;
      RECT 1845.815000 0.000000 1850.070000 0.630000 ;
      RECT 1841.310000 0.000000 1845.395000 0.630000 ;
      RECT 1836.720000 0.000000 1840.890000 0.630000 ;
      RECT 1832.045000 0.000000 1836.300000 0.630000 ;
      RECT 1827.710000 0.000000 1831.625000 0.630000 ;
      RECT 1822.950000 0.000000 1827.290000 0.630000 ;
      RECT 1818.700000 0.000000 1822.530000 0.630000 ;
      RECT 1814.110000 0.000000 1818.280000 0.630000 ;
      RECT 1809.520000 0.000000 1813.690000 0.630000 ;
      RECT 1805.015000 0.000000 1809.100000 0.630000 ;
      RECT 1800.425000 0.000000 1804.595000 0.630000 ;
      RECT 1795.835000 0.000000 1800.005000 0.630000 ;
      RECT 1791.330000 0.000000 1795.415000 0.630000 ;
      RECT 1786.740000 0.000000 1790.910000 0.630000 ;
      RECT 1782.150000 0.000000 1786.320000 0.630000 ;
      RECT 1777.645000 0.000000 1781.730000 0.630000 ;
      RECT 1773.140000 0.000000 1777.225000 0.630000 ;
      RECT 1768.635000 0.000000 1772.720000 0.630000 ;
      RECT 1764.045000 0.000000 1768.215000 0.630000 ;
      RECT 1759.625000 0.000000 1763.625000 0.630000 ;
      RECT 1755.035000 0.000000 1759.205000 0.630000 ;
      RECT 1750.530000 0.000000 1754.615000 0.630000 ;
      RECT 1745.940000 0.000000 1750.110000 0.630000 ;
      RECT 1741.435000 0.000000 1745.520000 0.630000 ;
      RECT 1736.760000 0.000000 1741.015000 0.630000 ;
      RECT 1732.425000 0.000000 1736.340000 0.630000 ;
      RECT 1727.665000 0.000000 1732.005000 0.630000 ;
      RECT 1723.245000 0.000000 1727.245000 0.630000 ;
      RECT 1718.655000 0.000000 1722.825000 0.630000 ;
      RECT 1714.065000 0.000000 1718.235000 0.630000 ;
      RECT 1709.560000 0.000000 1713.645000 0.630000 ;
      RECT 1704.970000 0.000000 1709.140000 0.630000 ;
      RECT 1700.465000 0.000000 1704.550000 0.630000 ;
      RECT 1695.960000 0.000000 1700.045000 0.630000 ;
      RECT 1691.370000 0.000000 1695.540000 0.630000 ;
      RECT 1686.865000 0.000000 1690.950000 0.630000 ;
      RECT 1682.275000 0.000000 1686.445000 0.630000 ;
      RECT 1677.685000 0.000000 1681.855000 0.630000 ;
      RECT 1673.265000 0.000000 1677.265000 0.630000 ;
      RECT 1668.675000 0.000000 1672.845000 0.630000 ;
      RECT 1664.085000 0.000000 1668.255000 0.630000 ;
      RECT 1659.580000 0.000000 1663.665000 0.630000 ;
      RECT 1654.905000 0.000000 1659.160000 0.630000 ;
      RECT 1650.485000 0.000000 1654.485000 0.630000 ;
      RECT 1645.810000 0.000000 1650.065000 0.630000 ;
      RECT 1641.390000 0.000000 1645.390000 0.630000 ;
      RECT 1636.800000 0.000000 1640.970000 0.630000 ;
      RECT 1632.295000 0.000000 1636.380000 0.630000 ;
      RECT 1627.620000 0.000000 1631.875000 0.630000 ;
      RECT 1623.200000 0.000000 1627.200000 0.630000 ;
      RECT 1618.525000 0.000000 1622.780000 0.630000 ;
      RECT 1614.190000 0.000000 1618.105000 0.630000 ;
      RECT 1609.515000 0.000000 1613.770000 0.630000 ;
      RECT 1605.010000 0.000000 1609.095000 0.630000 ;
      RECT 1600.420000 0.000000 1604.590000 0.630000 ;
      RECT 1595.830000 0.000000 1600.000000 0.630000 ;
      RECT 1591.325000 0.000000 1595.410000 0.630000 ;
      RECT 1586.735000 0.000000 1590.905000 0.630000 ;
      RECT 1582.230000 0.000000 1586.315000 0.630000 ;
      RECT 1577.725000 0.000000 1581.810000 0.630000 ;
      RECT 1573.135000 0.000000 1577.305000 0.630000 ;
      RECT 1568.545000 0.000000 1572.715000 0.630000 ;
      RECT 1564.125000 0.000000 1568.125000 0.630000 ;
      RECT 1559.450000 0.000000 1563.705000 0.630000 ;
      RECT 1555.030000 0.000000 1559.030000 0.630000 ;
      RECT 1550.440000 0.000000 1554.610000 0.630000 ;
      RECT 1545.850000 0.000000 1550.020000 0.630000 ;
      RECT 1541.345000 0.000000 1545.430000 0.630000 ;
      RECT 1536.670000 0.000000 1540.925000 0.630000 ;
      RECT 1532.165000 0.000000 1536.250000 0.630000 ;
      RECT 1527.575000 0.000000 1531.745000 0.630000 ;
      RECT 1523.155000 0.000000 1527.155000 0.630000 ;
      RECT 1518.565000 0.000000 1522.735000 0.630000 ;
      RECT 1514.060000 0.000000 1518.145000 0.630000 ;
      RECT 1509.385000 0.000000 1513.640000 0.630000 ;
      RECT 1505.050000 0.000000 1508.965000 0.630000 ;
      RECT 1500.290000 0.000000 1504.630000 0.630000 ;
      RECT 1495.955000 0.000000 1499.870000 0.630000 ;
      RECT 1491.280000 0.000000 1495.535000 0.630000 ;
      RECT 1486.775000 0.000000 1490.860000 0.630000 ;
      RECT 1482.185000 0.000000 1486.355000 0.630000 ;
      RECT 1477.595000 0.000000 1481.765000 0.630000 ;
      RECT 1473.005000 0.000000 1477.175000 0.630000 ;
      RECT 1468.500000 0.000000 1472.585000 0.630000 ;
      RECT 1463.995000 0.000000 1468.080000 0.630000 ;
      RECT 1459.490000 0.000000 1463.575000 0.630000 ;
      RECT 1454.900000 0.000000 1459.070000 0.630000 ;
      RECT 1450.310000 0.000000 1454.480000 0.630000 ;
      RECT 1445.890000 0.000000 1449.890000 0.630000 ;
      RECT 1441.215000 0.000000 1445.470000 0.630000 ;
      RECT 1436.710000 0.000000 1440.795000 0.630000 ;
      RECT 1432.205000 0.000000 1436.290000 0.630000 ;
      RECT 1427.615000 0.000000 1431.785000 0.630000 ;
      RECT 1423.110000 0.000000 1427.195000 0.630000 ;
      RECT 1418.435000 0.000000 1422.690000 0.630000 ;
      RECT 1413.930000 0.000000 1418.015000 0.630000 ;
      RECT 1409.340000 0.000000 1413.510000 0.630000 ;
      RECT 1404.920000 0.000000 1408.920000 0.630000 ;
      RECT 1400.245000 0.000000 1404.500000 0.630000 ;
      RECT 1395.825000 0.000000 1399.825000 0.630000 ;
      RECT 1391.150000 0.000000 1395.405000 0.630000 ;
      RECT 1386.815000 0.000000 1390.730000 0.630000 ;
      RECT 1382.055000 0.000000 1386.395000 0.630000 ;
      RECT 1377.635000 0.000000 1381.635000 0.630000 ;
      RECT 1373.045000 0.000000 1377.215000 0.630000 ;
      RECT 1368.540000 0.000000 1372.625000 0.630000 ;
      RECT 1363.950000 0.000000 1368.120000 0.630000 ;
      RECT 1359.360000 0.000000 1363.530000 0.630000 ;
      RECT 1354.770000 0.000000 1358.940000 0.630000 ;
      RECT 1350.265000 0.000000 1354.350000 0.630000 ;
      RECT 1345.760000 0.000000 1349.845000 0.630000 ;
      RECT 1341.170000 0.000000 1345.340000 0.630000 ;
      RECT 1336.665000 0.000000 1340.750000 0.630000 ;
      RECT 1332.075000 0.000000 1336.245000 0.630000 ;
      RECT 1327.655000 0.000000 1331.655000 0.630000 ;
      RECT 1323.065000 0.000000 1327.235000 0.630000 ;
      RECT 1318.475000 0.000000 1322.645000 0.630000 ;
      RECT 1313.970000 0.000000 1318.055000 0.630000 ;
      RECT 1309.380000 0.000000 1313.550000 0.630000 ;
      RECT 1304.790000 0.000000 1308.960000 0.630000 ;
      RECT 1300.200000 0.000000 1304.370000 0.630000 ;
      RECT 1295.695000 0.000000 1299.780000 0.630000 ;
      RECT 1291.105000 0.000000 1295.275000 0.630000 ;
      RECT 1286.685000 0.000000 1290.685000 0.630000 ;
      RECT 1282.010000 0.000000 1286.265000 0.630000 ;
      RECT 1277.590000 0.000000 1281.590000 0.630000 ;
      RECT 1272.915000 0.000000 1277.170000 0.630000 ;
      RECT 1268.580000 0.000000 1272.495000 0.630000 ;
      RECT 1263.905000 0.000000 1268.160000 0.630000 ;
      RECT 1259.400000 0.000000 1263.485000 0.630000 ;
      RECT 1254.810000 0.000000 1258.980000 0.630000 ;
      RECT 1250.305000 0.000000 1254.390000 0.630000 ;
      RECT 1245.630000 0.000000 1249.885000 0.630000 ;
      RECT 1241.125000 0.000000 1245.210000 0.630000 ;
      RECT 1236.535000 0.000000 1240.705000 0.630000 ;
      RECT 1232.030000 0.000000 1236.115000 0.630000 ;
      RECT 1227.525000 0.000000 1231.610000 0.630000 ;
      RECT 1222.935000 0.000000 1227.105000 0.630000 ;
      RECT 1218.515000 0.000000 1222.515000 0.630000 ;
      RECT 1213.840000 0.000000 1218.095000 0.630000 ;
      RECT 1209.250000 0.000000 1213.420000 0.630000 ;
      RECT 1204.830000 0.000000 1208.830000 0.630000 ;
      RECT 1200.240000 0.000000 1204.410000 0.630000 ;
      RECT 1195.735000 0.000000 1199.820000 0.630000 ;
      RECT 1191.145000 0.000000 1195.315000 0.630000 ;
      RECT 1186.640000 0.000000 1190.725000 0.630000 ;
      RECT 1182.050000 0.000000 1186.220000 0.630000 ;
      RECT 1177.545000 0.000000 1181.630000 0.630000 ;
      RECT 1172.870000 0.000000 1177.125000 0.630000 ;
      RECT 1168.620000 0.000000 1172.450000 0.630000 ;
      RECT 1163.860000 0.000000 1168.200000 0.630000 ;
      RECT 1159.525000 0.000000 1163.440000 0.630000 ;
      RECT 1154.850000 0.000000 1159.105000 0.630000 ;
      RECT 1150.345000 0.000000 1154.430000 0.630000 ;
      RECT 1145.755000 0.000000 1149.925000 0.630000 ;
      RECT 1141.250000 0.000000 1145.335000 0.630000 ;
      RECT 1136.660000 0.000000 1140.830000 0.630000 ;
      RECT 1132.155000 0.000000 1136.240000 0.630000 ;
      RECT 1127.480000 0.000000 1131.735000 0.630000 ;
      RECT 1122.975000 0.000000 1127.060000 0.630000 ;
      RECT 1118.385000 0.000000 1122.555000 0.630000 ;
      RECT 1113.795000 0.000000 1117.965000 0.630000 ;
      RECT 1109.460000 0.000000 1113.375000 0.630000 ;
      RECT 1104.785000 0.000000 1109.040000 0.630000 ;
      RECT 1100.365000 0.000000 1104.365000 0.630000 ;
      RECT 1095.775000 0.000000 1099.945000 0.630000 ;
      RECT 1091.185000 0.000000 1095.355000 0.630000 ;
      RECT 1086.680000 0.000000 1090.765000 0.630000 ;
      RECT 1082.090000 0.000000 1086.260000 0.630000 ;
      RECT 1077.500000 0.000000 1081.670000 0.630000 ;
      RECT 1072.995000 0.000000 1077.080000 0.630000 ;
      RECT 1068.405000 0.000000 1072.575000 0.630000 ;
      RECT 1063.815000 0.000000 1067.985000 0.630000 ;
      RECT 1059.310000 0.000000 1063.395000 0.630000 ;
      RECT 1054.635000 0.000000 1058.890000 0.630000 ;
      RECT 1050.385000 0.000000 1054.215000 0.630000 ;
      RECT 1045.710000 0.000000 1049.965000 0.630000 ;
      RECT 1041.290000 0.000000 1045.290000 0.630000 ;
      RECT 1036.615000 0.000000 1040.870000 0.630000 ;
      RECT 1032.110000 0.000000 1036.195000 0.630000 ;
      RECT 1027.520000 0.000000 1031.690000 0.630000 ;
      RECT 1023.015000 0.000000 1027.100000 0.630000 ;
      RECT 1018.340000 0.000000 1022.595000 0.630000 ;
      RECT 1013.920000 0.000000 1017.920000 0.630000 ;
      RECT 1009.245000 0.000000 1013.500000 0.630000 ;
      RECT 1004.740000 0.000000 1008.825000 0.630000 ;
      RECT 1000.150000 0.000000 1004.320000 0.630000 ;
      RECT 995.560000 0.000000 999.730000 0.630000 ;
      RECT 991.225000 0.000000 995.140000 0.630000 ;
      RECT 986.635000 0.000000 990.805000 0.630000 ;
      RECT 982.045000 0.000000 986.215000 0.630000 ;
      RECT 977.540000 0.000000 981.625000 0.630000 ;
      RECT 972.950000 0.000000 977.120000 0.630000 ;
      RECT 968.445000 0.000000 972.530000 0.630000 ;
      RECT 963.855000 0.000000 968.025000 0.630000 ;
      RECT 959.265000 0.000000 963.435000 0.630000 ;
      RECT 954.760000 0.000000 958.845000 0.630000 ;
      RECT 950.170000 0.000000 954.340000 0.630000 ;
      RECT 945.580000 0.000000 949.750000 0.630000 ;
      RECT 941.075000 0.000000 945.160000 0.630000 ;
      RECT 936.400000 0.000000 940.655000 0.630000 ;
      RECT 932.150000 0.000000 935.980000 0.630000 ;
      RECT 927.475000 0.000000 931.730000 0.630000 ;
      RECT 922.970000 0.000000 927.055000 0.630000 ;
      RECT 918.380000 0.000000 922.550000 0.630000 ;
      RECT 913.875000 0.000000 917.960000 0.630000 ;
      RECT 909.285000 0.000000 913.455000 0.630000 ;
      RECT 904.780000 0.000000 908.865000 0.630000 ;
      RECT 900.105000 0.000000 904.360000 0.630000 ;
      RECT 895.685000 0.000000 899.685000 0.630000 ;
      RECT 891.010000 0.000000 895.265000 0.630000 ;
      RECT 886.505000 0.000000 890.590000 0.630000 ;
      RECT 882.000000 0.000000 886.085000 0.630000 ;
      RECT 877.325000 0.000000 881.580000 0.630000 ;
      RECT 872.990000 0.000000 876.905000 0.630000 ;
      RECT 868.400000 0.000000 872.570000 0.630000 ;
      RECT 863.810000 0.000000 867.980000 0.630000 ;
      RECT 859.305000 0.000000 863.390000 0.630000 ;
      RECT 854.715000 0.000000 858.885000 0.630000 ;
      RECT 850.125000 0.000000 854.295000 0.630000 ;
      RECT 845.620000 0.000000 849.705000 0.630000 ;
      RECT 841.030000 0.000000 845.200000 0.630000 ;
      RECT 836.525000 0.000000 840.610000 0.630000 ;
      RECT 831.935000 0.000000 836.105000 0.630000 ;
      RECT 827.345000 0.000000 831.515000 0.630000 ;
      RECT 822.925000 0.000000 826.925000 0.630000 ;
      RECT 818.165000 0.000000 822.505000 0.630000 ;
      RECT 813.915000 0.000000 817.745000 0.630000 ;
      RECT 809.240000 0.000000 813.495000 0.630000 ;
      RECT 804.735000 0.000000 808.820000 0.630000 ;
      RECT 800.145000 0.000000 804.315000 0.630000 ;
      RECT 795.640000 0.000000 799.725000 0.630000 ;
      RECT 790.965000 0.000000 795.220000 0.630000 ;
      RECT 786.545000 0.000000 790.545000 0.630000 ;
      RECT 781.870000 0.000000 786.125000 0.630000 ;
      RECT 777.535000 0.000000 781.450000 0.630000 ;
      RECT 772.775000 0.000000 777.115000 0.630000 ;
      RECT 768.270000 0.000000 772.355000 0.630000 ;
      RECT 763.765000 0.000000 767.850000 0.630000 ;
      RECT 759.090000 0.000000 763.345000 0.630000 ;
      RECT 754.670000 0.000000 758.670000 0.630000 ;
      RECT 750.165000 0.000000 754.250000 0.630000 ;
      RECT 745.575000 0.000000 749.745000 0.630000 ;
      RECT 741.070000 0.000000 745.155000 0.630000 ;
      RECT 736.480000 0.000000 740.650000 0.630000 ;
      RECT 731.890000 0.000000 736.060000 0.630000 ;
      RECT 727.385000 0.000000 731.470000 0.630000 ;
      RECT 722.795000 0.000000 726.965000 0.630000 ;
      RECT 718.205000 0.000000 722.375000 0.630000 ;
      RECT 713.700000 0.000000 717.785000 0.630000 ;
      RECT 709.195000 0.000000 713.280000 0.630000 ;
      RECT 704.690000 0.000000 708.775000 0.630000 ;
      RECT 700.100000 0.000000 704.270000 0.630000 ;
      RECT 695.595000 0.000000 699.680000 0.630000 ;
      RECT 691.005000 0.000000 695.175000 0.630000 ;
      RECT 686.500000 0.000000 690.585000 0.630000 ;
      RECT 681.910000 0.000000 686.080000 0.630000 ;
      RECT 677.405000 0.000000 681.490000 0.630000 ;
      RECT 672.730000 0.000000 676.985000 0.630000 ;
      RECT 668.310000 0.000000 672.310000 0.630000 ;
      RECT 663.635000 0.000000 667.890000 0.630000 ;
      RECT 659.130000 0.000000 663.215000 0.630000 ;
      RECT 654.540000 0.000000 658.710000 0.630000 ;
      RECT 650.120000 0.000000 654.120000 0.630000 ;
      RECT 645.530000 0.000000 649.700000 0.630000 ;
      RECT 641.025000 0.000000 645.110000 0.630000 ;
      RECT 636.435000 0.000000 640.605000 0.630000 ;
      RECT 631.930000 0.000000 636.015000 0.630000 ;
      RECT 627.340000 0.000000 631.510000 0.630000 ;
      RECT 622.835000 0.000000 626.920000 0.630000 ;
      RECT 618.245000 0.000000 622.415000 0.630000 ;
      RECT 613.740000 0.000000 617.825000 0.630000 ;
      RECT 609.150000 0.000000 613.320000 0.630000 ;
      RECT 604.730000 0.000000 608.730000 0.630000 ;
      RECT 600.140000 0.000000 604.310000 0.630000 ;
      RECT 595.635000 0.000000 599.720000 0.630000 ;
      RECT 591.045000 0.000000 595.215000 0.630000 ;
      RECT 586.625000 0.000000 590.625000 0.630000 ;
      RECT 581.950000 0.000000 586.205000 0.630000 ;
      RECT 577.445000 0.000000 581.530000 0.630000 ;
      RECT 572.855000 0.000000 577.025000 0.630000 ;
      RECT 568.350000 0.000000 572.435000 0.630000 ;
      RECT 563.675000 0.000000 567.930000 0.630000 ;
      RECT 559.255000 0.000000 563.255000 0.630000 ;
      RECT 554.580000 0.000000 558.835000 0.630000 ;
      RECT 550.245000 0.000000 554.160000 0.630000 ;
      RECT 545.570000 0.000000 549.825000 0.630000 ;
      RECT 541.065000 0.000000 545.150000 0.630000 ;
      RECT 536.475000 0.000000 540.645000 0.630000 ;
      RECT 531.970000 0.000000 536.055000 0.630000 ;
      RECT 527.295000 0.000000 531.550000 0.630000 ;
      RECT 522.875000 0.000000 526.875000 0.630000 ;
      RECT 518.285000 0.000000 522.455000 0.630000 ;
      RECT 513.780000 0.000000 517.865000 0.630000 ;
      RECT 509.190000 0.000000 513.360000 0.630000 ;
      RECT 504.600000 0.000000 508.770000 0.630000 ;
      RECT 500.095000 0.000000 504.180000 0.630000 ;
      RECT 495.505000 0.000000 499.675000 0.630000 ;
      RECT 490.915000 0.000000 495.085000 0.630000 ;
      RECT 486.495000 0.000000 490.495000 0.630000 ;
      RECT 481.905000 0.000000 486.075000 0.630000 ;
      RECT 477.400000 0.000000 481.485000 0.630000 ;
      RECT 472.810000 0.000000 476.980000 0.630000 ;
      RECT 468.220000 0.000000 472.390000 0.630000 ;
      RECT 463.715000 0.000000 467.800000 0.630000 ;
      RECT 459.210000 0.000000 463.295000 0.630000 ;
      RECT 454.620000 0.000000 458.790000 0.630000 ;
      RECT 450.115000 0.000000 454.200000 0.630000 ;
      RECT 445.440000 0.000000 449.695000 0.630000 ;
      RECT 441.105000 0.000000 445.020000 0.630000 ;
      RECT 436.345000 0.000000 440.685000 0.630000 ;
      RECT 431.925000 0.000000 435.925000 0.630000 ;
      RECT 427.335000 0.000000 431.505000 0.630000 ;
      RECT 422.830000 0.000000 426.915000 0.630000 ;
      RECT 418.240000 0.000000 422.410000 0.630000 ;
      RECT 413.735000 0.000000 417.820000 0.630000 ;
      RECT 409.060000 0.000000 413.315000 0.630000 ;
      RECT 404.640000 0.000000 408.640000 0.630000 ;
      RECT 400.050000 0.000000 404.220000 0.630000 ;
      RECT 395.460000 0.000000 399.630000 0.630000 ;
      RECT 390.955000 0.000000 395.040000 0.630000 ;
      RECT 386.365000 0.000000 390.535000 0.630000 ;
      RECT 381.945000 0.000000 385.945000 0.630000 ;
      RECT 377.270000 0.000000 381.525000 0.630000 ;
      RECT 372.765000 0.000000 376.850000 0.630000 ;
      RECT 368.260000 0.000000 372.345000 0.630000 ;
      RECT 363.670000 0.000000 367.840000 0.630000 ;
      RECT 359.165000 0.000000 363.250000 0.630000 ;
      RECT 354.575000 0.000000 358.745000 0.630000 ;
      RECT 349.985000 0.000000 354.155000 0.630000 ;
      RECT 345.480000 0.000000 349.565000 0.630000 ;
      RECT 340.975000 0.000000 345.060000 0.630000 ;
      RECT 336.300000 0.000000 340.555000 0.630000 ;
      RECT 331.880000 0.000000 335.880000 0.630000 ;
      RECT 327.205000 0.000000 331.460000 0.630000 ;
      RECT 322.870000 0.000000 326.785000 0.630000 ;
      RECT 318.110000 0.000000 322.450000 0.630000 ;
      RECT 313.690000 0.000000 317.690000 0.630000 ;
      RECT 309.100000 0.000000 313.270000 0.630000 ;
      RECT 304.595000 0.000000 308.680000 0.630000 ;
      RECT 299.920000 0.000000 304.175000 0.630000 ;
      RECT 295.500000 0.000000 299.500000 0.630000 ;
      RECT 290.825000 0.000000 295.080000 0.630000 ;
      RECT 286.405000 0.000000 290.405000 0.630000 ;
      RECT 281.815000 0.000000 285.985000 0.630000 ;
      RECT 277.225000 0.000000 281.395000 0.630000 ;
      RECT 272.720000 0.000000 276.805000 0.630000 ;
      RECT 268.130000 0.000000 272.300000 0.630000 ;
      RECT 263.540000 0.000000 267.710000 0.630000 ;
      RECT 259.120000 0.000000 263.120000 0.630000 ;
      RECT 254.530000 0.000000 258.700000 0.630000 ;
      RECT 250.025000 0.000000 254.110000 0.630000 ;
      RECT 245.435000 0.000000 249.605000 0.630000 ;
      RECT 240.845000 0.000000 245.015000 0.630000 ;
      RECT 236.340000 0.000000 240.425000 0.630000 ;
      RECT 231.750000 0.000000 235.920000 0.630000 ;
      RECT 227.245000 0.000000 231.330000 0.630000 ;
      RECT 222.740000 0.000000 226.825000 0.630000 ;
      RECT 218.065000 0.000000 222.320000 0.630000 ;
      RECT 213.645000 0.000000 217.645000 0.630000 ;
      RECT 208.970000 0.000000 213.225000 0.630000 ;
      RECT 204.465000 0.000000 208.550000 0.630000 ;
      RECT 199.960000 0.000000 204.045000 0.630000 ;
      RECT 195.455000 0.000000 199.540000 0.630000 ;
      RECT 190.865000 0.000000 195.035000 0.630000 ;
      RECT 186.360000 0.000000 190.445000 0.630000 ;
      RECT 181.685000 0.000000 185.940000 0.630000 ;
      RECT 177.265000 0.000000 181.265000 0.630000 ;
      RECT 172.590000 0.000000 176.845000 0.630000 ;
      RECT 168.170000 0.000000 172.170000 0.630000 ;
      RECT 163.580000 0.000000 167.750000 0.630000 ;
      RECT 158.990000 0.000000 163.160000 0.630000 ;
      RECT 154.485000 0.000000 158.570000 0.630000 ;
      RECT 149.895000 0.000000 154.065000 0.630000 ;
      RECT 145.305000 0.000000 149.475000 0.630000 ;
      RECT 140.885000 0.000000 144.885000 0.630000 ;
      RECT 136.295000 0.000000 140.465000 0.630000 ;
      RECT 131.790000 0.000000 135.875000 0.630000 ;
      RECT 127.200000 0.000000 131.370000 0.630000 ;
      RECT 122.610000 0.000000 126.780000 0.630000 ;
      RECT 118.105000 0.000000 122.190000 0.630000 ;
      RECT 113.515000 0.000000 117.685000 0.630000 ;
      RECT 109.010000 0.000000 113.095000 0.630000 ;
      RECT 104.505000 0.000000 108.590000 0.630000 ;
      RECT 99.830000 0.000000 104.085000 0.630000 ;
      RECT 95.495000 0.000000 99.410000 0.630000 ;
      RECT 90.735000 0.000000 95.075000 0.630000 ;
      RECT 86.315000 0.000000 90.315000 0.630000 ;
      RECT 81.725000 0.000000 85.895000 0.630000 ;
      RECT 77.220000 0.000000 81.305000 0.630000 ;
      RECT 72.545000 0.000000 76.800000 0.630000 ;
      RECT 68.125000 0.000000 72.125000 0.630000 ;
      RECT 63.450000 0.000000 67.705000 0.630000 ;
      RECT 59.030000 0.000000 63.030000 0.630000 ;
      RECT 54.355000 0.000000 58.610000 0.630000 ;
      RECT 49.935000 0.000000 53.935000 0.630000 ;
      RECT 45.345000 0.000000 49.515000 0.630000 ;
      RECT 40.840000 0.000000 44.925000 0.630000 ;
      RECT 36.335000 0.000000 40.420000 0.630000 ;
      RECT 31.830000 0.000000 35.915000 0.630000 ;
      RECT 27.240000 0.000000 31.410000 0.630000 ;
      RECT 22.735000 0.000000 26.820000 0.630000 ;
      RECT 18.145000 0.000000 22.315000 0.630000 ;
      RECT 13.555000 0.000000 17.725000 0.630000 ;
      RECT 9.050000 0.000000 13.135000 0.630000 ;
      RECT 4.460000 0.000000 8.630000 0.630000 ;
      RECT 2.505000 0.000000 4.040000 0.625000 ;
      RECT 0.000000 0.000000 2.085000 0.625000 ;
    LAYER met3 ;
      RECT 0.000000 2176.750000 2300.000000 2219.180000 ;
      RECT 0.000000 2176.350000 2298.900000 2176.750000 ;
      RECT 1.100000 2175.850000 2298.900000 2176.350000 ;
      RECT 1.100000 2175.450000 2300.000000 2175.850000 ;
      RECT 0.000000 2137.250000 2300.000000 2175.450000 ;
      RECT 1.100000 2136.550000 2300.000000 2137.250000 ;
      RECT 1.100000 2136.350000 2298.900000 2136.550000 ;
      RECT 0.000000 2135.650000 2298.900000 2136.350000 ;
      RECT 0.000000 2096.250000 2300.000000 2135.650000 ;
      RECT 1.100000 2095.350000 2300.000000 2096.250000 ;
      RECT 0.000000 2094.650000 2300.000000 2095.350000 ;
      RECT 0.000000 2093.750000 2298.900000 2094.650000 ;
      RECT 0.000000 2055.050000 2300.000000 2093.750000 ;
      RECT 1.100000 2054.150000 2300.000000 2055.050000 ;
      RECT 0.000000 2052.750000 2300.000000 2054.150000 ;
      RECT 0.000000 2051.850000 2298.900000 2052.750000 ;
      RECT 0.000000 2013.950000 2300.000000 2051.850000 ;
      RECT 1.100000 2013.050000 2300.000000 2013.950000 ;
      RECT 0.000000 2010.850000 2300.000000 2013.050000 ;
      RECT 0.000000 2009.950000 2298.900000 2010.850000 ;
      RECT 0.000000 1972.950000 2300.000000 2009.950000 ;
      RECT 1.100000 1972.050000 2300.000000 1972.950000 ;
      RECT 0.000000 1969.050000 2300.000000 1972.050000 ;
      RECT 0.000000 1968.150000 2298.900000 1969.050000 ;
      RECT 0.000000 1931.750000 2300.000000 1968.150000 ;
      RECT 1.100000 1930.850000 2300.000000 1931.750000 ;
      RECT 0.000000 1927.050000 2300.000000 1930.850000 ;
      RECT 0.000000 1926.150000 2298.900000 1927.050000 ;
      RECT 0.000000 1890.750000 2300.000000 1926.150000 ;
      RECT 1.100000 1889.850000 2300.000000 1890.750000 ;
      RECT 0.000000 1885.150000 2300.000000 1889.850000 ;
      RECT 0.000000 1884.250000 2298.900000 1885.150000 ;
      RECT 0.000000 1849.650000 2300.000000 1884.250000 ;
      RECT 1.100000 1848.750000 2300.000000 1849.650000 ;
      RECT 0.000000 1843.350000 2300.000000 1848.750000 ;
      RECT 0.000000 1842.450000 2298.900000 1843.350000 ;
      RECT 0.000000 1808.550000 2300.000000 1842.450000 ;
      RECT 1.100000 1807.650000 2300.000000 1808.550000 ;
      RECT 0.000000 1801.350000 2300.000000 1807.650000 ;
      RECT 0.000000 1800.450000 2298.900000 1801.350000 ;
      RECT 0.000000 1767.450000 2300.000000 1800.450000 ;
      RECT 1.100000 1766.550000 2300.000000 1767.450000 ;
      RECT 0.000000 1759.550000 2300.000000 1766.550000 ;
      RECT 0.000000 1758.650000 2298.900000 1759.550000 ;
      RECT 0.000000 1726.350000 2300.000000 1758.650000 ;
      RECT 1.100000 1725.450000 2300.000000 1726.350000 ;
      RECT 0.000000 1717.650000 2300.000000 1725.450000 ;
      RECT 0.000000 1716.750000 2298.900000 1717.650000 ;
      RECT 0.000000 1685.150000 2300.000000 1716.750000 ;
      RECT 1.100000 1684.250000 2300.000000 1685.150000 ;
      RECT 0.000000 1675.750000 2300.000000 1684.250000 ;
      RECT 0.000000 1674.850000 2298.900000 1675.750000 ;
      RECT 0.000000 1644.150000 2300.000000 1674.850000 ;
      RECT 1.100000 1643.250000 2300.000000 1644.150000 ;
      RECT 0.000000 1633.850000 2300.000000 1643.250000 ;
      RECT 0.000000 1632.950000 2298.900000 1633.850000 ;
      RECT 0.000000 1603.050000 2300.000000 1632.950000 ;
      RECT 1.100000 1602.150000 2300.000000 1603.050000 ;
      RECT 0.000000 1591.950000 2300.000000 1602.150000 ;
      RECT 0.000000 1591.050000 2298.900000 1591.950000 ;
      RECT 0.000000 1561.950000 2300.000000 1591.050000 ;
      RECT 1.100000 1561.050000 2300.000000 1561.950000 ;
      RECT 0.000000 1550.050000 2300.000000 1561.050000 ;
      RECT 0.000000 1549.150000 2298.900000 1550.050000 ;
      RECT 0.000000 1520.950000 2300.000000 1549.150000 ;
      RECT 1.100000 1520.050000 2300.000000 1520.950000 ;
      RECT 0.000000 1508.150000 2300.000000 1520.050000 ;
      RECT 0.000000 1507.250000 2298.900000 1508.150000 ;
      RECT 0.000000 1479.750000 2300.000000 1507.250000 ;
      RECT 1.100000 1478.850000 2300.000000 1479.750000 ;
      RECT 0.000000 1466.350000 2300.000000 1478.850000 ;
      RECT 0.000000 1465.450000 2298.900000 1466.350000 ;
      RECT 0.000000 1438.650000 2300.000000 1465.450000 ;
      RECT 1.100000 1437.750000 2300.000000 1438.650000 ;
      RECT 0.000000 1424.350000 2300.000000 1437.750000 ;
      RECT 0.000000 1423.450000 2298.900000 1424.350000 ;
      RECT 0.000000 1397.550000 2300.000000 1423.450000 ;
      RECT 1.100000 1396.650000 2300.000000 1397.550000 ;
      RECT 0.000000 1382.550000 2300.000000 1396.650000 ;
      RECT 0.000000 1381.650000 2298.900000 1382.550000 ;
      RECT 0.000000 1356.450000 2300.000000 1381.650000 ;
      RECT 1.100000 1355.550000 2300.000000 1356.450000 ;
      RECT 0.000000 1340.650000 2300.000000 1355.550000 ;
      RECT 0.000000 1339.750000 2298.900000 1340.650000 ;
      RECT 0.000000 1315.350000 2300.000000 1339.750000 ;
      RECT 1.100000 1314.450000 2300.000000 1315.350000 ;
      RECT 0.000000 1298.750000 2300.000000 1314.450000 ;
      RECT 0.000000 1297.850000 2298.900000 1298.750000 ;
      RECT 0.000000 1274.350000 2300.000000 1297.850000 ;
      RECT 1.100000 1273.450000 2300.000000 1274.350000 ;
      RECT 0.000000 1256.950000 2300.000000 1273.450000 ;
      RECT 0.000000 1256.050000 2298.900000 1256.950000 ;
      RECT 0.000000 1233.150000 2300.000000 1256.050000 ;
      RECT 1.100000 1232.250000 2300.000000 1233.150000 ;
      RECT 0.000000 1214.950000 2300.000000 1232.250000 ;
      RECT 0.000000 1214.050000 2298.900000 1214.950000 ;
      RECT 0.000000 1192.150000 2300.000000 1214.050000 ;
      RECT 1.100000 1191.250000 2300.000000 1192.150000 ;
      RECT 0.000000 1173.150000 2300.000000 1191.250000 ;
      RECT 0.000000 1172.250000 2298.900000 1173.150000 ;
      RECT 0.000000 1151.050000 2300.000000 1172.250000 ;
      RECT 1.100000 1150.150000 2300.000000 1151.050000 ;
      RECT 0.000000 1131.250000 2300.000000 1150.150000 ;
      RECT 0.000000 1130.350000 2298.900000 1131.250000 ;
      RECT 0.000000 1109.850000 2300.000000 1130.350000 ;
      RECT 1.100000 1108.950000 2300.000000 1109.850000 ;
      RECT 0.000000 1089.350000 2300.000000 1108.950000 ;
      RECT 0.000000 1088.450000 2298.900000 1089.350000 ;
      RECT 0.000000 1068.850000 2300.000000 1088.450000 ;
      RECT 1.100000 1067.950000 2300.000000 1068.850000 ;
      RECT 0.000000 1047.550000 2300.000000 1067.950000 ;
      RECT 0.000000 1046.650000 2298.900000 1047.550000 ;
      RECT 0.000000 1027.750000 2300.000000 1046.650000 ;
      RECT 1.100000 1026.850000 2300.000000 1027.750000 ;
      RECT 0.000000 1005.550000 2300.000000 1026.850000 ;
      RECT 0.000000 1004.650000 2298.900000 1005.550000 ;
      RECT 0.000000 986.550000 2300.000000 1004.650000 ;
      RECT 1.100000 985.650000 2300.000000 986.550000 ;
      RECT 0.000000 963.750000 2300.000000 985.650000 ;
      RECT 0.000000 962.850000 2298.900000 963.750000 ;
      RECT 0.000000 945.550000 2300.000000 962.850000 ;
      RECT 1.100000 944.650000 2300.000000 945.550000 ;
      RECT 0.000000 921.850000 2300.000000 944.650000 ;
      RECT 0.000000 920.950000 2298.900000 921.850000 ;
      RECT 0.000000 904.450000 2300.000000 920.950000 ;
      RECT 1.100000 903.550000 2300.000000 904.450000 ;
      RECT 0.000000 879.950000 2300.000000 903.550000 ;
      RECT 0.000000 879.050000 2298.900000 879.950000 ;
      RECT 0.000000 863.350000 2300.000000 879.050000 ;
      RECT 1.100000 862.450000 2300.000000 863.350000 ;
      RECT 0.000000 838.050000 2300.000000 862.450000 ;
      RECT 0.000000 837.150000 2298.900000 838.050000 ;
      RECT 0.000000 822.250000 2300.000000 837.150000 ;
      RECT 1.100000 821.350000 2300.000000 822.250000 ;
      RECT 0.000000 796.150000 2300.000000 821.350000 ;
      RECT 0.000000 795.250000 2298.900000 796.150000 ;
      RECT 0.000000 781.050000 2300.000000 795.250000 ;
      RECT 1.100000 780.150000 2300.000000 781.050000 ;
      RECT 0.000000 754.250000 2300.000000 780.150000 ;
      RECT 0.000000 753.350000 2298.900000 754.250000 ;
      RECT 0.000000 740.050000 2300.000000 753.350000 ;
      RECT 1.100000 739.150000 2300.000000 740.050000 ;
      RECT 0.000000 712.350000 2300.000000 739.150000 ;
      RECT 0.000000 711.450000 2298.900000 712.350000 ;
      RECT 0.000000 698.950000 2300.000000 711.450000 ;
      RECT 1.100000 698.050000 2300.000000 698.950000 ;
      RECT 0.000000 670.550000 2300.000000 698.050000 ;
      RECT 0.000000 669.650000 2298.900000 670.550000 ;
      RECT 0.000000 657.850000 2300.000000 669.650000 ;
      RECT 1.100000 656.950000 2300.000000 657.850000 ;
      RECT 0.000000 628.550000 2300.000000 656.950000 ;
      RECT 0.000000 627.650000 2298.900000 628.550000 ;
      RECT 0.000000 616.750000 2300.000000 627.650000 ;
      RECT 1.100000 615.850000 2300.000000 616.750000 ;
      RECT 0.000000 586.750000 2300.000000 615.850000 ;
      RECT 0.000000 585.850000 2298.900000 586.750000 ;
      RECT 0.000000 575.750000 2300.000000 585.850000 ;
      RECT 1.100000 574.850000 2300.000000 575.750000 ;
      RECT 0.000000 544.850000 2300.000000 574.850000 ;
      RECT 0.000000 543.950000 2298.900000 544.850000 ;
      RECT 0.000000 534.550000 2300.000000 543.950000 ;
      RECT 1.100000 533.650000 2300.000000 534.550000 ;
      RECT 0.000000 502.950000 2300.000000 533.650000 ;
      RECT 0.000000 502.050000 2298.900000 502.950000 ;
      RECT 0.000000 493.450000 2300.000000 502.050000 ;
      RECT 1.100000 492.550000 2300.000000 493.450000 ;
      RECT 0.000000 461.050000 2300.000000 492.550000 ;
      RECT 0.000000 460.150000 2298.900000 461.050000 ;
      RECT 0.000000 452.350000 2300.000000 460.150000 ;
      RECT 1.100000 451.450000 2300.000000 452.350000 ;
      RECT 0.000000 419.150000 2300.000000 451.450000 ;
      RECT 0.000000 418.250000 2298.900000 419.150000 ;
      RECT 0.000000 411.250000 2300.000000 418.250000 ;
      RECT 1.100000 410.350000 2300.000000 411.250000 ;
      RECT 0.000000 377.250000 2300.000000 410.350000 ;
      RECT 0.000000 376.350000 2298.900000 377.250000 ;
      RECT 0.000000 370.150000 2300.000000 376.350000 ;
      RECT 1.100000 369.250000 2300.000000 370.150000 ;
      RECT 0.000000 335.350000 2300.000000 369.250000 ;
      RECT 0.000000 334.450000 2298.900000 335.350000 ;
      RECT 0.000000 329.050000 2300.000000 334.450000 ;
      RECT 1.100000 328.150000 2300.000000 329.050000 ;
      RECT 0.000000 293.550000 2300.000000 328.150000 ;
      RECT 0.000000 292.650000 2298.900000 293.550000 ;
      RECT 0.000000 288.050000 2300.000000 292.650000 ;
      RECT 1.100000 287.150000 2300.000000 288.050000 ;
      RECT 0.000000 251.550000 2300.000000 287.150000 ;
      RECT 0.000000 250.650000 2298.900000 251.550000 ;
      RECT 0.000000 246.950000 2300.000000 250.650000 ;
      RECT 1.100000 246.050000 2300.000000 246.950000 ;
      RECT 0.000000 209.750000 2300.000000 246.050000 ;
      RECT 0.000000 208.850000 2298.900000 209.750000 ;
      RECT 0.000000 205.750000 2300.000000 208.850000 ;
      RECT 1.100000 204.850000 2300.000000 205.750000 ;
      RECT 0.000000 167.850000 2300.000000 204.850000 ;
      RECT 0.000000 166.950000 2298.900000 167.850000 ;
      RECT 0.000000 164.650000 2300.000000 166.950000 ;
      RECT 1.100000 163.750000 2300.000000 164.650000 ;
      RECT 0.000000 125.950000 2300.000000 163.750000 ;
      RECT 0.000000 125.050000 2298.900000 125.950000 ;
      RECT 0.000000 123.650000 2300.000000 125.050000 ;
      RECT 1.100000 122.750000 2300.000000 123.650000 ;
      RECT 0.000000 84.150000 2300.000000 122.750000 ;
      RECT 0.000000 83.250000 2298.900000 84.150000 ;
      RECT 0.000000 58.020000 2300.000000 83.250000 ;
      RECT 1.100000 57.120000 2300.000000 58.020000 ;
      RECT 0.000000 42.250000 2300.000000 57.120000 ;
      RECT 0.000000 41.450000 2298.900000 42.250000 ;
      RECT 1.100000 41.350000 2298.900000 41.450000 ;
      RECT 1.100000 40.550000 2300.000000 41.350000 ;
      RECT 0.000000 4.550000 2300.000000 40.550000 ;
      RECT 0.000000 3.650000 2298.900000 4.550000 ;
      RECT 0.000000 2.750000 2300.000000 3.650000 ;
      RECT 1.100000 1.850000 2300.000000 2.750000 ;
      RECT 0.000000 0.000000 2300.000000 1.850000 ;
    LAYER met4 ;
      RECT 0.000000 2197.360000 2300.000000 2219.180000 ;
      RECT 35.200000 2177.360000 2264.340000 2197.360000 ;
      RECT 2260.140000 39.440000 2264.340000 2177.360000 ;
      RECT 55.200000 39.440000 2244.340000 2177.360000 ;
      RECT 35.200000 39.440000 39.400000 2177.360000 ;
      RECT 2280.140000 19.440000 2300.000000 2197.360000 ;
      RECT 35.200000 19.440000 2264.340000 39.440000 ;
      RECT 0.000000 19.440000 19.400000 2197.360000 ;
      RECT 0.000000 0.000000 2300.000000 19.440000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
